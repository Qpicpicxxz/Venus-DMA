# Confidential Information of ARM, Inc.
# Use subject to ARM license.
# Copyright (c) 2024 ARM, Inc.

# ACI Version r1p1

# Reifier 4.0.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;

#name: High Density Dual Port SRAM RVT RVT Compiler | LOGIC0040LL 40nm Process 0.589um^2 Bit Cell
#version: r1p1
#comment: 
#configuration:  -activity_factor 50 -back_biasing off -bits 64 -bmux on -bus_notation on -check_instname on -diodes on -drive 6 -ema on -frequency 1.0 -instname SRAMdpw64d256 -left_bus_delim "[" -mux 4 -mvt "" -name_case upper -power_type otc -prefix "" -pwr_gnd_rename vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -retention on -right_bus_delim "]" -rows_p_bl 256 -ser none -site_def off -top_layer m5-m10 -words 256 -write_mask off -write_thru off -corners ff_1p21v_1p21v_0c,ff_1p21v_1p21v_125c,ff_1p21v_1p21v_m40c,ss_0p99v_0p99v_0c,ss_0p99v_0p99v_125c,ss_0p99v_0p99v_m40c,tt_1p10v_1p10v_125c,tt_1p10v_1p10v_25c,tt_1p10v_1p10v_85c
MACRO SRAMdpw64d256
  FOREIGN SRAMdpw64d256 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 442.43 BY 69.945 ;
  CLASS BLOCK ;
  PIN RET1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 221.955 0.0 222.095 0.25 ;
      LAYER M2 ;
      RECT 221.955 0.0 222.095 0.25 ;
      LAYER M1 ;
      RECT 221.955 0.0 222.095 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END RET1N
  PIN COLLDISN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 229.855 0.0 229.995 0.25 ;
      LAYER M2 ;
      RECT 229.855 0.0 229.995 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END COLLDISN
  PIN SOA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 211.51 0.0 211.65 0.25 ;
      LAYER M3 ;
      RECT 211.51 0.0 211.65 0.25 ;
      LAYER M2 ;
      RECT 211.51 0.0 211.65 0.25 ;
      LAYER M1 ;
      RECT 211.51 0.0 211.65 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END SOA[0]
  PIN SOA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 230.6 0.0 230.74 0.25 ;
      LAYER M2 ;
      RECT 230.6 0.0 230.74 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END SOA[1]
  PIN CLKA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 211.21 0.0 211.35 0.25 ;
      LAYER M2 ;
      RECT 211.21 0.0 211.35 0.25 ;
      LAYER M1 ;
      RECT 211.21 0.0 211.35 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CLKA
  PIN CLKB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 231.02 0.0 231.16 0.25 ;
      LAYER M2 ;
      RECT 231.02 0.0 231.16 0.25 ;
      LAYER M3 ;
      RECT 231.02 0.0 231.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CLKB
  PIN SOB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 210.605 0.0 210.745 0.25 ;
      LAYER M3 ;
      RECT 210.605 0.0 210.745 0.25 ;
      LAYER M2 ;
      RECT 210.605 0.0 210.745 0.25 ;
      LAYER M1 ;
      RECT 210.605 0.0 210.745 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END SOB[0]
  PIN SOB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 231.685 0.0 231.825 0.25 ;
      LAYER M2 ;
      RECT 231.685 0.0 231.825 0.25 ;
      LAYER M3 ;
      RECT 231.685 0.0 231.825 0.25 ;
      LAYER M4 ;
      RECT 231.685 0.0 231.825 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END SOB[1]
  PIN EMAWA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 207.03 0.0 207.17 0.25 ;
      LAYER M2 ;
      RECT 207.03 0.0 207.17 0.25 ;
      LAYER M1 ;
      RECT 207.03 0.0 207.17 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAWA[0]
  PIN EMAWB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 235.235 0.0 235.375 0.25 ;
      LAYER M2 ;
      RECT 235.235 0.0 235.375 0.25 ;
      LAYER M3 ;
      RECT 235.235 0.0 235.375 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAWB[0]
  PIN AYA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 206.29 0.0 206.43 0.25 ;
      LAYER M2 ;
      RECT 206.29 0.0 206.43 0.25 ;
      LAYER M1 ;
      RECT 206.29 0.0 206.43 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[0]
  PIN AYB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 235.68 0.0 235.82 0.25 ;
      LAYER M2 ;
      RECT 235.68 0.0 235.82 0.25 ;
      LAYER M3 ;
      RECT 235.68 0.0 235.82 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[0]
  PIN TAA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 205.565 0.0 205.705 0.25 ;
      LAYER M2 ;
      RECT 205.565 0.0 205.705 0.25 ;
      LAYER M1 ;
      RECT 205.565 0.0 205.705 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[0]
  PIN TAB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 237.36 0.0 237.5 0.25 ;
      LAYER M2 ;
      RECT 237.36 0.0 237.5 0.25 ;
      LAYER M3 ;
      RECT 237.36 0.0 237.5 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[0]
  PIN AA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 205.26 0.0 205.4 0.25 ;
      LAYER M2 ;
      RECT 205.26 0.0 205.4 0.25 ;
      LAYER M1 ;
      RECT 205.26 0.0 205.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[0]
  PIN AB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 237.77 0.0 237.91 0.25 ;
      LAYER M2 ;
      RECT 237.77 0.0 237.91 0.25 ;
      LAYER M3 ;
      RECT 237.77 0.0 237.91 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[0]
  PIN EMAWA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 203.02 0.0 203.16 0.25 ;
      LAYER M2 ;
      RECT 203.02 0.0 203.16 0.25 ;
      LAYER M1 ;
      RECT 203.02 0.0 203.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAWA[1]
  PIN EMAWB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 239.27 0.0 239.41 0.25 ;
      LAYER M2 ;
      RECT 239.27 0.0 239.41 0.25 ;
      LAYER M3 ;
      RECT 239.27 0.0 239.41 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAWB[1]
  PIN EMAA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 202.64 0.0 202.78 0.25 ;
      LAYER M2 ;
      RECT 202.64 0.0 202.78 0.25 ;
      LAYER M1 ;
      RECT 202.64 0.0 202.78 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAA[0]
  PIN EMAB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 239.65 0.0 239.79 0.25 ;
      LAYER M2 ;
      RECT 239.65 0.0 239.79 0.25 ;
      LAYER M3 ;
      RECT 239.65 0.0 239.79 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAB[0]
  PIN AYA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 201.825 0.0 201.965 0.25 ;
      LAYER M2 ;
      RECT 201.825 0.0 201.965 0.25 ;
      LAYER M1 ;
      RECT 201.825 0.0 201.965 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[1]
  PIN AYB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 240.27 0.0 240.41 0.25 ;
      LAYER M2 ;
      RECT 240.27 0.0 240.41 0.25 ;
      LAYER M3 ;
      RECT 240.27 0.0 240.41 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[1]
  PIN TAA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 201.225 0.0 201.365 0.25 ;
      LAYER M2 ;
      RECT 201.225 0.0 201.365 0.25 ;
      LAYER M1 ;
      RECT 201.225 0.0 201.365 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[1]
  PIN TAB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 240.705 0.0 240.845 0.25 ;
      LAYER M2 ;
      RECT 240.705 0.0 240.845 0.25 ;
      LAYER M3 ;
      RECT 240.705 0.0 240.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[1]
  PIN AA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 200.775 0.0 200.915 0.25 ;
      LAYER M2 ;
      RECT 200.775 0.0 200.915 0.25 ;
      LAYER M1 ;
      RECT 200.775 0.0 200.915 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[1]
  PIN AB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 241.26 0.0 241.4 0.25 ;
      LAYER M2 ;
      RECT 241.26 0.0 241.4 0.25 ;
      LAYER M3 ;
      RECT 241.26 0.0 241.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[1]
  PIN EMAA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 199.8 0.0 199.94 0.25 ;
      LAYER M2 ;
      RECT 199.8 0.0 199.94 0.25 ;
      LAYER M1 ;
      RECT 199.8 0.0 199.94 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAA[2]
  PIN EMAB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 242.705 0.0 242.845 0.25 ;
      LAYER M2 ;
      RECT 242.705 0.0 242.845 0.25 ;
      LAYER M3 ;
      RECT 242.705 0.0 242.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAB[2]
  PIN TDB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 199.185 0.0 199.325 0.25 ;
      LAYER M2 ;
      RECT 199.185 0.0 199.325 0.25 ;
      LAYER M1 ;
      RECT 199.185 0.0 199.325 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[31]
  PIN TDB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 243.065 0.0 243.205 0.25 ;
      LAYER M2 ;
      RECT 243.065 0.0 243.205 0.25 ;
      LAYER M3 ;
      RECT 243.065 0.0 243.205 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[32]
  PIN EMAA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 198.905 0.0 199.045 0.25 ;
      LAYER M2 ;
      RECT 198.905 0.0 199.045 0.25 ;
      LAYER M1 ;
      RECT 198.905 0.0 199.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAA[1]
  PIN EMAB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 243.385 0.0 243.525 0.25 ;
      LAYER M2 ;
      RECT 243.385 0.0 243.525 0.25 ;
      LAYER M3 ;
      RECT 243.385 0.0 243.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAB[1]
  PIN QB[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 198.625 0.0 198.765 0.25 ;
      LAYER M3 ;
      RECT 198.625 0.0 198.765 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[31]
  PIN QB[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 243.665 0.0 243.805 0.25 ;
      LAYER M4 ;
      RECT 243.665 0.0 243.805 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[32]
  PIN DB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 198.275 0.0 198.415 0.25 ;
      LAYER M2 ;
      RECT 198.275 0.0 198.415 0.25 ;
      LAYER M1 ;
      RECT 198.275 0.0 198.415 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[31]
  PIN DB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 244.035 0.0 244.175 0.25 ;
      LAYER M2 ;
      RECT 244.035 0.0 244.175 0.25 ;
      LAYER M3 ;
      RECT 244.035 0.0 244.175 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[32]
  PIN DA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 194.545 0.0 194.685 0.25 ;
      LAYER M3 ;
      RECT 194.545 0.0 194.685 0.25 ;
      LAYER M2 ;
      RECT 194.545 0.0 194.685 0.25 ;
      LAYER M1 ;
      RECT 194.545 0.0 194.685 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[31]
  PIN DA[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 247.745 0.0 247.885 0.25 ;
      LAYER M2 ;
      RECT 247.745 0.0 247.885 0.25 ;
      LAYER M3 ;
      RECT 247.745 0.0 247.885 0.25 ;
      LAYER M4 ;
      RECT 247.745 0.0 247.885 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[32]
  PIN QA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 194.245 0.0 194.385 0.25 ;
      LAYER M3 ;
      RECT 194.245 0.0 194.385 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[31]
  PIN QA[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 248.135 0.0 248.275 0.25 ;
      LAYER M4 ;
      RECT 248.135 0.0 248.275 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[32]
  PIN TDA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 193.685 0.0 193.825 0.25 ;
      LAYER M2 ;
      RECT 193.685 0.0 193.825 0.25 ;
      LAYER M1 ;
      RECT 193.685 0.0 193.825 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[31]
  PIN TDA[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 248.815 0.0 248.955 0.25 ;
      LAYER M2 ;
      RECT 248.815 0.0 248.955 0.25 ;
      LAYER M3 ;
      RECT 248.815 0.0 248.955 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[32]
  PIN TDB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 193.125 0.0 193.265 0.25 ;
      LAYER M2 ;
      RECT 193.125 0.0 193.265 0.25 ;
      LAYER M1 ;
      RECT 193.125 0.0 193.265 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[30]
  PIN TDB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 249.38 0.0 249.52 0.25 ;
      LAYER M2 ;
      RECT 249.38 0.0 249.52 0.25 ;
      LAYER M3 ;
      RECT 249.38 0.0 249.52 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[33]
  PIN QB[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 192.425 0.0 192.565 0.25 ;
      LAYER M3 ;
      RECT 192.425 0.0 192.565 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[30]
  PIN QB[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 250.0 0.0 250.14 0.25 ;
      LAYER M4 ;
      RECT 250.0 0.0 250.14 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[33]
  PIN DB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 192.035 0.0 192.175 0.25 ;
      LAYER M3 ;
      RECT 192.035 0.0 192.175 0.25 ;
      LAYER M2 ;
      RECT 192.035 0.0 192.175 0.25 ;
      LAYER M1 ;
      RECT 192.035 0.0 192.175 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[30]
  PIN DB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 250.295 0.0 250.435 0.25 ;
      LAYER M2 ;
      RECT 250.295 0.0 250.435 0.25 ;
      LAYER M3 ;
      RECT 250.295 0.0 250.435 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[33]
  PIN SEA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 190.505 0.0 190.645 0.25 ;
      LAYER M2 ;
      RECT 190.505 0.0 190.645 0.25 ;
      LAYER M1 ;
      RECT 190.505 0.0 190.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END SEA
  PIN SEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 251.52 0.0 251.66 0.25 ;
      LAYER M2 ;
      RECT 251.52 0.0 251.66 0.25 ;
      LAYER M3 ;
      RECT 251.52 0.0 251.66 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END SEB
  PIN AYA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 190.13 0.0 190.27 0.25 ;
      LAYER M2 ;
      RECT 190.13 0.0 190.27 0.25 ;
      LAYER M1 ;
      RECT 190.13 0.0 190.27 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[2]
  PIN AYB[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 251.82 0.0 251.96 0.25 ;
      LAYER M2 ;
      RECT 251.82 0.0 251.96 0.25 ;
      LAYER M3 ;
      RECT 251.82 0.0 251.96 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[2]
  PIN TAA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 189.825 0.0 189.965 0.25 ;
      LAYER M2 ;
      RECT 189.825 0.0 189.965 0.25 ;
      LAYER M1 ;
      RECT 189.825 0.0 189.965 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[2]
  PIN TAB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 252.585 0.0 252.725 0.25 ;
      LAYER M2 ;
      RECT 252.585 0.0 252.725 0.25 ;
      LAYER M3 ;
      RECT 252.585 0.0 252.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[2]
  PIN AA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 189.53 0.0 189.67 0.25 ;
      LAYER M2 ;
      RECT 189.53 0.0 189.67 0.25 ;
      LAYER M1 ;
      RECT 189.53 0.0 189.67 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[2]
  PIN AB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 252.88 0.0 253.02 0.25 ;
      LAYER M2 ;
      RECT 252.88 0.0 253.02 0.25 ;
      LAYER M3 ;
      RECT 252.88 0.0 253.02 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[2]
  PIN DA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 188.345 0.0 188.485 0.25 ;
      LAYER M3 ;
      RECT 188.345 0.0 188.485 0.25 ;
      LAYER M2 ;
      RECT 188.345 0.0 188.485 0.25 ;
      LAYER M1 ;
      RECT 188.345 0.0 188.485 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[30]
  PIN DA[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 253.945 0.0 254.085 0.25 ;
      LAYER M2 ;
      RECT 253.945 0.0 254.085 0.25 ;
      LAYER M3 ;
      RECT 253.945 0.0 254.085 0.25 ;
      LAYER M4 ;
      RECT 253.945 0.0 254.085 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[33]
  PIN QA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 187.955 0.0 188.095 0.25 ;
      LAYER M3 ;
      RECT 187.955 0.0 188.095 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[30]
  PIN QA[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 254.335 0.0 254.475 0.25 ;
      LAYER M4 ;
      RECT 254.335 0.0 254.475 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[33]
  PIN TDA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 187.34 0.0 187.48 0.25 ;
      LAYER M2 ;
      RECT 187.34 0.0 187.48 0.25 ;
      LAYER M1 ;
      RECT 187.34 0.0 187.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[30]
  PIN TDA[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 254.935 0.0 255.075 0.25 ;
      LAYER M2 ;
      RECT 254.935 0.0 255.075 0.25 ;
      LAYER M3 ;
      RECT 254.935 0.0 255.075 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[33]
  PIN TDB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 186.9 0.0 187.04 0.25 ;
      LAYER M2 ;
      RECT 186.9 0.0 187.04 0.25 ;
      LAYER M1 ;
      RECT 186.9 0.0 187.04 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[29]
  PIN TDB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 255.505 0.0 255.645 0.25 ;
      LAYER M2 ;
      RECT 255.505 0.0 255.645 0.25 ;
      LAYER M3 ;
      RECT 255.505 0.0 255.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[34]
  PIN AYA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 186.585 0.0 186.725 0.25 ;
      LAYER M2 ;
      RECT 186.585 0.0 186.725 0.25 ;
      LAYER M1 ;
      RECT 186.585 0.0 186.725 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[3]
  PIN AYB[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 255.785 0.0 255.925 0.25 ;
      LAYER M2 ;
      RECT 255.785 0.0 255.925 0.25 ;
      LAYER M3 ;
      RECT 255.785 0.0 255.925 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[3]
  PIN QB[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 186.225 0.0 186.365 0.25 ;
      LAYER M3 ;
      RECT 186.225 0.0 186.365 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[29]
  PIN QB[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 256.065 0.0 256.205 0.25 ;
      LAYER M4 ;
      RECT 256.065 0.0 256.205 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[34]
  PIN DB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 185.92 0.0 186.06 0.25 ;
      LAYER M3 ;
      RECT 185.92 0.0 186.06 0.25 ;
      LAYER M2 ;
      RECT 185.92 0.0 186.06 0.25 ;
      LAYER M1 ;
      RECT 185.92 0.0 186.06 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[29]
  PIN DB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 256.455 0.0 256.595 0.25 ;
      LAYER M2 ;
      RECT 256.455 0.0 256.595 0.25 ;
      LAYER M3 ;
      RECT 256.455 0.0 256.595 0.25 ;
      LAYER M4 ;
      RECT 256.455 0.0 256.595 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[34]
  PIN TAA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 185.64 0.0 185.78 0.25 ;
      LAYER M2 ;
      RECT 185.64 0.0 185.78 0.25 ;
      LAYER M1 ;
      RECT 185.64 0.0 185.78 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[3]
  PIN TAB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 256.745 0.0 256.885 0.25 ;
      LAYER M2 ;
      RECT 256.745 0.0 256.885 0.25 ;
      LAYER M3 ;
      RECT 256.745 0.0 256.885 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[3]
  PIN AA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 184.63 0.0 184.77 0.25 ;
      LAYER M2 ;
      RECT 184.63 0.0 184.77 0.25 ;
      LAYER M1 ;
      RECT 184.63 0.0 184.77 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[3]
  PIN AB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 257.595 0.0 257.735 0.25 ;
      LAYER M2 ;
      RECT 257.595 0.0 257.735 0.25 ;
      LAYER M3 ;
      RECT 257.595 0.0 257.735 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[3]
  PIN AYA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 182.38 0.0 182.52 0.25 ;
      LAYER M2 ;
      RECT 182.38 0.0 182.52 0.25 ;
      LAYER M1 ;
      RECT 182.38 0.0 182.52 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[4]
  PIN AYB[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 259.845 0.0 259.985 0.25 ;
      LAYER M2 ;
      RECT 259.845 0.0 259.985 0.25 ;
      LAYER M3 ;
      RECT 259.845 0.0 259.985 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[4]
  PIN DA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 182.1 0.0 182.24 0.25 ;
      LAYER M3 ;
      RECT 182.1 0.0 182.24 0.25 ;
      LAYER M2 ;
      RECT 182.1 0.0 182.24 0.25 ;
      LAYER M1 ;
      RECT 182.1 0.0 182.24 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[29]
  PIN DA[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 260.145 0.0 260.285 0.25 ;
      LAYER M2 ;
      RECT 260.145 0.0 260.285 0.25 ;
      LAYER M3 ;
      RECT 260.145 0.0 260.285 0.25 ;
      LAYER M4 ;
      RECT 260.145 0.0 260.285 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[34]
  PIN QA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 181.755 0.0 181.895 0.25 ;
      LAYER M3 ;
      RECT 181.755 0.0 181.895 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[29]
  PIN QA[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 260.535 0.0 260.675 0.25 ;
      LAYER M4 ;
      RECT 260.535 0.0 260.675 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[34]
  PIN TAA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 181.435 0.0 181.575 0.25 ;
      LAYER M2 ;
      RECT 181.435 0.0 181.575 0.25 ;
      LAYER M1 ;
      RECT 181.435 0.0 181.575 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[4]
  PIN TAB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 260.84 0.0 260.98 0.25 ;
      LAYER M2 ;
      RECT 260.84 0.0 260.98 0.25 ;
      LAYER M3 ;
      RECT 260.84 0.0 260.98 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[4]
  PIN TDA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 181.105 0.0 181.245 0.25 ;
      LAYER M2 ;
      RECT 181.105 0.0 181.245 0.25 ;
      LAYER M1 ;
      RECT 181.105 0.0 181.245 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[29]
  PIN TDA[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 261.135 0.0 261.275 0.25 ;
      LAYER M2 ;
      RECT 261.135 0.0 261.275 0.25 ;
      LAYER M3 ;
      RECT 261.135 0.0 261.275 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[34]
  PIN AA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 180.82 0.0 180.96 0.25 ;
      LAYER M2 ;
      RECT 180.82 0.0 180.96 0.25 ;
      LAYER M1 ;
      RECT 180.82 0.0 180.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[4]
  PIN AB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 261.455 0.0 261.595 0.25 ;
      LAYER M2 ;
      RECT 261.455 0.0 261.595 0.25 ;
      LAYER M3 ;
      RECT 261.455 0.0 261.595 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[4]
  PIN TDB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 180.54 0.0 180.68 0.25 ;
      LAYER M2 ;
      RECT 180.54 0.0 180.68 0.25 ;
      LAYER M1 ;
      RECT 180.54 0.0 180.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[28]
  PIN TDB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 261.735 0.0 261.875 0.25 ;
      LAYER M2 ;
      RECT 261.735 0.0 261.875 0.25 ;
      LAYER M3 ;
      RECT 261.735 0.0 261.875 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[35]
  PIN DFTRAMBYP
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 180.26 0.0 180.4 0.25 ;
      LAYER M2 ;
      RECT 180.26 0.0 180.4 0.25 ;
      LAYER M1 ;
      RECT 180.26 0.0 180.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DFTRAMBYP
  PIN QB[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 262.265 0.0 262.405 0.25 ;
      LAYER M4 ;
      RECT 262.265 0.0 262.405 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[35]
  PIN QB[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 179.98 0.0 180.12 0.25 ;
      LAYER M3 ;
      RECT 179.98 0.0 180.12 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[28]
  PIN TENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 262.545 0.0 262.685 0.25 ;
      LAYER M2 ;
      RECT 262.545 0.0 262.685 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TENB
  PIN TENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 179.585 0.0 179.725 0.25 ;
      LAYER M1 ;
      RECT 179.585 0.0 179.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TENA
  PIN DB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 262.825 0.0 262.965 0.25 ;
      LAYER M2 ;
      RECT 262.825 0.0 262.965 0.25 ;
      LAYER M3 ;
      RECT 262.825 0.0 262.965 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[35]
  PIN DB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 179.275 0.0 179.415 0.25 ;
      LAYER M2 ;
      RECT 179.275 0.0 179.415 0.25 ;
      LAYER M1 ;
      RECT 179.275 0.0 179.415 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[28]
  PIN DA[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 266.345 0.0 266.485 0.25 ;
      LAYER M2 ;
      RECT 266.345 0.0 266.485 0.25 ;
      LAYER M3 ;
      RECT 266.345 0.0 266.485 0.25 ;
      LAYER M4 ;
      RECT 266.345 0.0 266.485 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[35]
  PIN DA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 175.945 0.0 176.085 0.25 ;
      LAYER M3 ;
      RECT 175.945 0.0 176.085 0.25 ;
      LAYER M2 ;
      RECT 175.945 0.0 176.085 0.25 ;
      LAYER M1 ;
      RECT 175.945 0.0 176.085 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[28]
  PIN QA[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 266.66 0.0 266.8 0.25 ;
      LAYER M4 ;
      RECT 266.66 0.0 266.8 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[35]
  PIN QA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 175.645 0.0 175.785 0.25 ;
      LAYER M3 ;
      RECT 175.645 0.0 175.785 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[28]
  PIN AYB[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 266.95 0.0 267.09 0.25 ;
      LAYER M2 ;
      RECT 266.95 0.0 267.09 0.25 ;
      LAYER M3 ;
      RECT 266.95 0.0 267.09 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[5]
  PIN AYA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 175.365 0.0 175.505 0.25 ;
      LAYER M2 ;
      RECT 175.365 0.0 175.505 0.25 ;
      LAYER M1 ;
      RECT 175.365 0.0 175.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[5]
  PIN TDA[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 267.23 0.0 267.37 0.25 ;
      LAYER M2 ;
      RECT 267.23 0.0 267.37 0.25 ;
      LAYER M3 ;
      RECT 267.23 0.0 267.37 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[35]
  PIN TDA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 175.065 0.0 175.205 0.25 ;
      LAYER M2 ;
      RECT 175.065 0.0 175.205 0.25 ;
      LAYER M1 ;
      RECT 175.065 0.0 175.205 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[28]
  PIN TAB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 267.51 0.0 267.65 0.25 ;
      LAYER M2 ;
      RECT 267.51 0.0 267.65 0.25 ;
      LAYER M3 ;
      RECT 267.51 0.0 267.65 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[5]
  PIN TAA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 174.78 0.0 174.92 0.25 ;
      LAYER M2 ;
      RECT 174.78 0.0 174.92 0.25 ;
      LAYER M1 ;
      RECT 174.78 0.0 174.92 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[5]
  PIN TDB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 267.795 0.0 267.935 0.25 ;
      LAYER M2 ;
      RECT 267.795 0.0 267.935 0.25 ;
      LAYER M3 ;
      RECT 267.795 0.0 267.935 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[36]
  PIN TDB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 174.5 0.0 174.64 0.25 ;
      LAYER M2 ;
      RECT 174.5 0.0 174.64 0.25 ;
      LAYER M1 ;
      RECT 174.5 0.0 174.64 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[27]
  PIN AB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 268.075 0.0 268.215 0.25 ;
      LAYER M2 ;
      RECT 268.075 0.0 268.215 0.25 ;
      LAYER M3 ;
      RECT 268.075 0.0 268.215 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[5]
  PIN AA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 174.175 0.0 174.315 0.25 ;
      LAYER M2 ;
      RECT 174.175 0.0 174.315 0.25 ;
      LAYER M1 ;
      RECT 174.175 0.0 174.315 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[5]
  PIN QB[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 268.465 0.0 268.605 0.25 ;
      LAYER M4 ;
      RECT 268.465 0.0 268.605 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[36]
  PIN QB[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 173.825 0.0 173.965 0.25 ;
      LAYER M3 ;
      RECT 173.825 0.0 173.965 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[27]
  PIN DB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 268.855 0.0 268.995 0.25 ;
      LAYER M2 ;
      RECT 268.855 0.0 268.995 0.25 ;
      LAYER M3 ;
      RECT 268.855 0.0 268.995 0.25 ;
      LAYER M4 ;
      RECT 268.855 0.0 268.995 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[36]
  PIN DB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 173.435 0.0 173.575 0.25 ;
      LAYER M3 ;
      RECT 173.435 0.0 173.575 0.25 ;
      LAYER M2 ;
      RECT 173.435 0.0 173.575 0.25 ;
      LAYER M1 ;
      RECT 173.435 0.0 173.575 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[27]
  PIN AYB[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 270.355 0.0 270.495 0.25 ;
      LAYER M2 ;
      RECT 270.355 0.0 270.495 0.25 ;
      LAYER M3 ;
      RECT 270.355 0.0 270.495 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[6]
  PIN AYA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 171.71 0.0 171.85 0.25 ;
      LAYER M2 ;
      RECT 171.71 0.0 171.85 0.25 ;
      LAYER M1 ;
      RECT 171.71 0.0 171.85 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[6]
  PIN TAB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 271.045 0.0 271.185 0.25 ;
      LAYER M2 ;
      RECT 271.045 0.0 271.185 0.25 ;
      LAYER M3 ;
      RECT 271.045 0.0 271.185 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[6]
  PIN TAA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 171.165 0.0 171.305 0.25 ;
      LAYER M2 ;
      RECT 171.165 0.0 171.305 0.25 ;
      LAYER M1 ;
      RECT 171.165 0.0 171.305 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[6]
  PIN AB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 271.325 0.0 271.465 0.25 ;
      LAYER M2 ;
      RECT 271.325 0.0 271.465 0.25 ;
      LAYER M3 ;
      RECT 271.325 0.0 271.465 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[6]
  PIN AA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 170.865 0.0 171.005 0.25 ;
      LAYER M2 ;
      RECT 170.865 0.0 171.005 0.25 ;
      LAYER M1 ;
      RECT 170.865 0.0 171.005 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[6]
  PIN DA[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 272.545 0.0 272.685 0.25 ;
      LAYER M2 ;
      RECT 272.545 0.0 272.685 0.25 ;
      LAYER M3 ;
      RECT 272.545 0.0 272.685 0.25 ;
      LAYER M4 ;
      RECT 272.545 0.0 272.685 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[36]
  PIN DA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 169.745 0.0 169.885 0.25 ;
      LAYER M3 ;
      RECT 169.745 0.0 169.885 0.25 ;
      LAYER M2 ;
      RECT 169.745 0.0 169.885 0.25 ;
      LAYER M1 ;
      RECT 169.745 0.0 169.885 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[27]
  PIN QA[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 272.935 0.0 273.075 0.25 ;
      LAYER M4 ;
      RECT 272.935 0.0 273.075 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[36]
  PIN QA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 169.355 0.0 169.495 0.25 ;
      LAYER M3 ;
      RECT 169.355 0.0 169.495 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[27]
  PIN TDA[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 273.52 0.0 273.66 0.25 ;
      LAYER M2 ;
      RECT 273.52 0.0 273.66 0.25 ;
      LAYER M3 ;
      RECT 273.52 0.0 273.66 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[36]
  PIN TDA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 168.795 0.0 168.935 0.25 ;
      LAYER M2 ;
      RECT 168.795 0.0 168.935 0.25 ;
      LAYER M1 ;
      RECT 168.795 0.0 168.935 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[27]
  PIN TDB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 274.09 0.0 274.23 0.25 ;
      LAYER M2 ;
      RECT 274.09 0.0 274.23 0.25 ;
      LAYER M3 ;
      RECT 274.09 0.0 274.23 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[37]
  PIN TDB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 168.225 0.0 168.365 0.25 ;
      LAYER M2 ;
      RECT 168.225 0.0 168.365 0.25 ;
      LAYER M1 ;
      RECT 168.225 0.0 168.365 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[26]
  PIN AYB[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 274.37 0.0 274.51 0.25 ;
      LAYER M2 ;
      RECT 274.37 0.0 274.51 0.25 ;
      LAYER M3 ;
      RECT 274.37 0.0 274.51 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYB[7]
  PIN AYA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 167.89 0.0 168.03 0.25 ;
      LAYER M2 ;
      RECT 167.89 0.0 168.03 0.25 ;
      LAYER M1 ;
      RECT 167.89 0.0 168.03 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END AYA[7]
  PIN QB[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 274.665 0.0 274.805 0.25 ;
      LAYER M4 ;
      RECT 274.665 0.0 274.805 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[37]
  PIN QB[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 167.585 0.0 167.725 0.25 ;
      LAYER M3 ;
      RECT 167.585 0.0 167.725 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[26]
  PIN TAB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 275.035 0.0 275.175 0.25 ;
      LAYER M2 ;
      RECT 275.035 0.0 275.175 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAB[7]
  PIN TAA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 167.285 0.0 167.425 0.25 ;
      LAYER M1 ;
      RECT 167.285 0.0 167.425 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TAA[7]
  PIN DB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 275.315 0.0 275.455 0.25 ;
      LAYER M2 ;
      RECT 275.315 0.0 275.455 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[37]
  PIN DB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 166.975 0.0 167.115 0.25 ;
      LAYER M2 ;
      RECT 166.975 0.0 167.115 0.25 ;
      LAYER M1 ;
      RECT 166.975 0.0 167.115 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[26]
  PIN AB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 276.385 0.0 276.525 0.25 ;
      LAYER M2 ;
      RECT 276.385 0.0 276.525 0.25 ;
      LAYER M3 ;
      RECT 276.385 0.0 276.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[7]
  PIN AA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 165.935 0.0 166.075 0.25 ;
      LAYER M2 ;
      RECT 165.935 0.0 166.075 0.25 ;
      LAYER M1 ;
      RECT 165.935 0.0 166.075 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[7]
  PIN DA[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 278.785 0.0 278.925 0.25 ;
      LAYER M2 ;
      RECT 278.785 0.0 278.925 0.25 ;
      LAYER M3 ;
      RECT 278.785 0.0 278.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[37]
  PIN DA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 163.495 0.0 163.635 0.25 ;
      LAYER M2 ;
      RECT 163.495 0.0 163.635 0.25 ;
      LAYER M1 ;
      RECT 163.495 0.0 163.635 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[26]
  PIN QA[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 279.135 0.0 279.275 0.25 ;
      LAYER M4 ;
      RECT 279.135 0.0 279.275 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[37]
  PIN QA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 163.185 0.0 163.325 0.25 ;
      LAYER M3 ;
      RECT 163.185 0.0 163.325 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[26]
  PIN TDA[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 279.845 0.0 279.985 0.25 ;
      LAYER M2 ;
      RECT 279.845 0.0 279.985 0.25 ;
      LAYER M3 ;
      RECT 279.845 0.0 279.985 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[37]
  PIN TDA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 162.615 0.0 162.755 0.25 ;
      LAYER M2 ;
      RECT 162.615 0.0 162.755 0.25 ;
      LAYER M1 ;
      RECT 162.615 0.0 162.755 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[26]
  PIN TDB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 280.41 0.0 280.55 0.25 ;
      LAYER M2 ;
      RECT 280.41 0.0 280.55 0.25 ;
      LAYER M3 ;
      RECT 280.41 0.0 280.55 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[38]
  PIN TDB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 162.025 0.0 162.165 0.25 ;
      LAYER M2 ;
      RECT 162.025 0.0 162.165 0.25 ;
      LAYER M1 ;
      RECT 162.025 0.0 162.165 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[25]
  PIN QB[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 280.865 0.0 281.005 0.25 ;
      LAYER M4 ;
      RECT 280.865 0.0 281.005 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[38]
  PIN QB[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 161.425 0.0 161.565 0.25 ;
      LAYER M3 ;
      RECT 161.425 0.0 161.565 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[25]
  PIN DB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 281.255 0.0 281.395 0.25 ;
      LAYER M2 ;
      RECT 281.255 0.0 281.395 0.25 ;
      LAYER M3 ;
      RECT 281.255 0.0 281.395 0.25 ;
      LAYER M4 ;
      RECT 281.255 0.0 281.395 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[38]
  PIN DB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 161.035 0.0 161.175 0.25 ;
      LAYER M3 ;
      RECT 161.035 0.0 161.175 0.25 ;
      LAYER M2 ;
      RECT 161.035 0.0 161.175 0.25 ;
      LAYER M1 ;
      RECT 161.035 0.0 161.175 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[25]
  PIN DA[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 284.945 0.0 285.085 0.25 ;
      LAYER M2 ;
      RECT 284.945 0.0 285.085 0.25 ;
      LAYER M3 ;
      RECT 284.945 0.0 285.085 0.25 ;
      LAYER M4 ;
      RECT 284.945 0.0 285.085 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[38]
  PIN DA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 157.345 0.0 157.485 0.25 ;
      LAYER M3 ;
      RECT 157.345 0.0 157.485 0.25 ;
      LAYER M2 ;
      RECT 157.345 0.0 157.485 0.25 ;
      LAYER M1 ;
      RECT 157.345 0.0 157.485 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[25]
  PIN QA[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 285.335 0.0 285.475 0.25 ;
      LAYER M4 ;
      RECT 285.335 0.0 285.475 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[38]
  PIN QA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 156.955 0.0 157.095 0.25 ;
      LAYER M3 ;
      RECT 156.955 0.0 157.095 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[25]
  PIN TDA[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 285.935 0.0 286.075 0.25 ;
      LAYER M2 ;
      RECT 285.935 0.0 286.075 0.25 ;
      LAYER M3 ;
      RECT 285.935 0.0 286.075 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[38]
  PIN TDA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 156.575 0.0 156.715 0.25 ;
      LAYER M2 ;
      RECT 156.575 0.0 156.715 0.25 ;
      LAYER M1 ;
      RECT 156.575 0.0 156.715 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[25]
  PIN TDB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 286.495 0.0 286.635 0.25 ;
      LAYER M2 ;
      RECT 286.495 0.0 286.635 0.25 ;
      LAYER M3 ;
      RECT 286.495 0.0 286.635 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[39]
  PIN TDB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 155.995 0.0 156.135 0.25 ;
      LAYER M2 ;
      RECT 155.995 0.0 156.135 0.25 ;
      LAYER M1 ;
      RECT 155.995 0.0 156.135 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[24]
  PIN QB[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 287.065 0.0 287.205 0.25 ;
      LAYER M4 ;
      RECT 287.065 0.0 287.205 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[39]
  PIN QB[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 155.06 0.0 155.2 0.25 ;
      LAYER M3 ;
      RECT 155.06 0.0 155.2 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[24]
  PIN DB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 287.625 0.0 287.765 0.25 ;
      LAYER M2 ;
      RECT 287.625 0.0 287.765 0.25 ;
      LAYER M3 ;
      RECT 287.625 0.0 287.765 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[39]
  PIN DB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 154.76 0.0 154.9 0.25 ;
      LAYER M1 ;
      RECT 154.76 0.0 154.9 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[24]
  PIN TCENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 288.575 0.0 288.715 0.25 ;
      LAYER M2 ;
      RECT 288.575 0.0 288.715 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TCENB
  PIN TCENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 153.825 0.0 153.965 0.25 ;
      LAYER M1 ;
      RECT 153.825 0.0 153.965 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TCENA
  PIN CENYB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 288.92 0.0 289.06 0.25 ;
      LAYER M2 ;
      RECT 288.92 0.0 289.06 0.25 ;
      LAYER M3 ;
      RECT 288.92 0.0 289.06 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END CENYB
  PIN CENYA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 153.515 0.0 153.655 0.25 ;
      LAYER M2 ;
      RECT 153.515 0.0 153.655 0.25 ;
      LAYER M1 ;
      RECT 153.515 0.0 153.655 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END CENYA
  PIN CENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 289.205 0.0 289.345 0.25 ;
      LAYER M2 ;
      RECT 289.205 0.0 289.345 0.25 ;
      LAYER M3 ;
      RECT 289.205 0.0 289.345 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CENB
  PIN CENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 153.14 0.0 153.28 0.25 ;
      LAYER M2 ;
      RECT 153.14 0.0 153.28 0.25 ;
      LAYER M1 ;
      RECT 153.14 0.0 153.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CENA
  PIN WENYB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 289.99 0.0 290.13 0.25 ;
      LAYER M2 ;
      RECT 289.99 0.0 290.13 0.25 ;
      LAYER M3 ;
      RECT 289.99 0.0 290.13 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END WENYB
  PIN WENYA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 152.37 0.0 152.51 0.25 ;
      LAYER M2 ;
      RECT 152.37 0.0 152.51 0.25 ;
      LAYER M1 ;
      RECT 152.37 0.0 152.51 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END WENYA
  PIN DA[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 290.905 0.0 291.045 0.25 ;
      LAYER M2 ;
      RECT 290.905 0.0 291.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[39]
  PIN DA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 151.44 0.0 151.58 0.25 ;
      LAYER M2 ;
      RECT 151.44 0.0 151.58 0.25 ;
      LAYER M1 ;
      RECT 151.44 0.0 151.58 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[24]
  PIN TWENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 291.25 0.0 291.39 0.25 ;
      LAYER M2 ;
      RECT 291.25 0.0 291.39 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TWENB
  PIN TWENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
      RECT 151.13 0.0 151.27 0.25 ;
      LAYER M1 ;
      RECT 151.13 0.0 151.27 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TWENA
  PIN QA[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 291.535 0.0 291.675 0.25 ;
      LAYER M4 ;
      RECT 291.535 0.0 291.675 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[39]
  PIN QA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 150.755 0.0 150.895 0.25 ;
      LAYER M3 ;
      RECT 150.755 0.0 150.895 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[24]
  PIN WENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 291.935 0.0 292.075 0.25 ;
      LAYER M2 ;
      RECT 291.935 0.0 292.075 0.25 ;
      LAYER M3 ;
      RECT 291.935 0.0 292.075 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END WENB
  PIN WENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 150.455 0.0 150.595 0.25 ;
      LAYER M2 ;
      RECT 150.455 0.0 150.595 0.25 ;
      LAYER M1 ;
      RECT 150.455 0.0 150.595 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END WENA
  PIN TDA[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 292.215 0.0 292.355 0.25 ;
      LAYER M2 ;
      RECT 292.215 0.0 292.355 0.25 ;
      LAYER M3 ;
      RECT 292.215 0.0 292.355 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[39]
  PIN TDA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 150.175 0.0 150.315 0.25 ;
      LAYER M2 ;
      RECT 150.175 0.0 150.315 0.25 ;
      LAYER M1 ;
      RECT 150.175 0.0 150.315 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[24]
  PIN TDB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 292.67 0.0 292.81 0.25 ;
      LAYER M2 ;
      RECT 292.67 0.0 292.81 0.25 ;
      LAYER M3 ;
      RECT 292.67 0.0 292.81 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[40]
  PIN TDB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 149.62 0.0 149.76 0.25 ;
      LAYER M2 ;
      RECT 149.62 0.0 149.76 0.25 ;
      LAYER M1 ;
      RECT 149.62 0.0 149.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[23]
  PIN QB[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 293.055 0.0 293.195 0.25 ;
      LAYER M2 ;
      RECT 293.055 0.0 293.195 0.25 ;
      LAYER M3 ;
      RECT 293.055 0.0 293.195 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[40]
  PIN QB[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 149.235 0.0 149.375 0.25 ;
      LAYER M2 ;
      RECT 149.235 0.0 149.375 0.25 ;
      LAYER M1 ;
      RECT 149.235 0.0 149.375 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[23]
  PIN DB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 293.83 0.0 293.97 0.25 ;
      LAYER M2 ;
      RECT 293.83 0.0 293.97 0.25 ;
      LAYER M3 ;
      RECT 293.83 0.0 293.97 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[40]
  PIN DB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 148.46 0.0 148.6 0.25 ;
      LAYER M2 ;
      RECT 148.46 0.0 148.6 0.25 ;
      LAYER M1 ;
      RECT 148.46 0.0 148.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[23]
  PIN DA[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 297.14 0.0 297.28 0.25 ;
      LAYER M2 ;
      RECT 297.14 0.0 297.28 0.25 ;
      LAYER M3 ;
      RECT 297.14 0.0 297.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[40]
  PIN DA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 145.15 0.0 145.29 0.25 ;
      LAYER M2 ;
      RECT 145.15 0.0 145.29 0.25 ;
      LAYER M1 ;
      RECT 145.15 0.0 145.29 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[23]
  PIN QA[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 297.925 0.0 298.065 0.25 ;
      LAYER M2 ;
      RECT 297.925 0.0 298.065 0.25 ;
      LAYER M3 ;
      RECT 297.925 0.0 298.065 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[40]
  PIN QA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 144.365 0.0 144.505 0.25 ;
      LAYER M2 ;
      RECT 144.365 0.0 144.505 0.25 ;
      LAYER M1 ;
      RECT 144.365 0.0 144.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[23]
  PIN TDA[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 298.305 0.0 298.445 0.25 ;
      LAYER M2 ;
      RECT 298.305 0.0 298.445 0.25 ;
      LAYER M3 ;
      RECT 298.305 0.0 298.445 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[40]
  PIN TDA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 143.985 0.0 144.125 0.25 ;
      LAYER M2 ;
      RECT 143.985 0.0 144.125 0.25 ;
      LAYER M1 ;
      RECT 143.985 0.0 144.125 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[23]
  PIN TDB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 298.87 0.0 299.01 0.25 ;
      LAYER M2 ;
      RECT 298.87 0.0 299.01 0.25 ;
      LAYER M3 ;
      RECT 298.87 0.0 299.01 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[41]
  PIN TDB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 143.42 0.0 143.56 0.25 ;
      LAYER M2 ;
      RECT 143.42 0.0 143.56 0.25 ;
      LAYER M1 ;
      RECT 143.42 0.0 143.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[22]
  PIN QB[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 299.255 0.0 299.395 0.25 ;
      LAYER M2 ;
      RECT 299.255 0.0 299.395 0.25 ;
      LAYER M3 ;
      RECT 299.255 0.0 299.395 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[41]
  PIN QB[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 143.035 0.0 143.175 0.25 ;
      LAYER M2 ;
      RECT 143.035 0.0 143.175 0.25 ;
      LAYER M1 ;
      RECT 143.035 0.0 143.175 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[22]
  PIN DB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 300.03 0.0 300.17 0.25 ;
      LAYER M2 ;
      RECT 300.03 0.0 300.17 0.25 ;
      LAYER M3 ;
      RECT 300.03 0.0 300.17 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[41]
  PIN DB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 142.26 0.0 142.4 0.25 ;
      LAYER M2 ;
      RECT 142.26 0.0 142.4 0.25 ;
      LAYER M1 ;
      RECT 142.26 0.0 142.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[22]
  PIN DA[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 303.34 0.0 303.48 0.25 ;
      LAYER M2 ;
      RECT 303.34 0.0 303.48 0.25 ;
      LAYER M3 ;
      RECT 303.34 0.0 303.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[41]
  PIN DA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 138.95 0.0 139.09 0.25 ;
      LAYER M2 ;
      RECT 138.95 0.0 139.09 0.25 ;
      LAYER M1 ;
      RECT 138.95 0.0 139.09 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[22]
  PIN QA[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 304.125 0.0 304.265 0.25 ;
      LAYER M2 ;
      RECT 304.125 0.0 304.265 0.25 ;
      LAYER M3 ;
      RECT 304.125 0.0 304.265 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[41]
  PIN QA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 138.165 0.0 138.305 0.25 ;
      LAYER M2 ;
      RECT 138.165 0.0 138.305 0.25 ;
      LAYER M1 ;
      RECT 138.165 0.0 138.305 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[22]
  PIN TDA[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 304.505 0.0 304.645 0.25 ;
      LAYER M2 ;
      RECT 304.505 0.0 304.645 0.25 ;
      LAYER M3 ;
      RECT 304.505 0.0 304.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[41]
  PIN TDA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 137.785 0.0 137.925 0.25 ;
      LAYER M2 ;
      RECT 137.785 0.0 137.925 0.25 ;
      LAYER M1 ;
      RECT 137.785 0.0 137.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[22]
  PIN TDB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 305.07 0.0 305.21 0.25 ;
      LAYER M2 ;
      RECT 305.07 0.0 305.21 0.25 ;
      LAYER M3 ;
      RECT 305.07 0.0 305.21 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[42]
  PIN TDB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 137.22 0.0 137.36 0.25 ;
      LAYER M2 ;
      RECT 137.22 0.0 137.36 0.25 ;
      LAYER M1 ;
      RECT 137.22 0.0 137.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[21]
  PIN QB[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 305.455 0.0 305.595 0.25 ;
      LAYER M2 ;
      RECT 305.455 0.0 305.595 0.25 ;
      LAYER M3 ;
      RECT 305.455 0.0 305.595 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[42]
  PIN QB[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 136.835 0.0 136.975 0.25 ;
      LAYER M2 ;
      RECT 136.835 0.0 136.975 0.25 ;
      LAYER M1 ;
      RECT 136.835 0.0 136.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[21]
  PIN DB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 306.23 0.0 306.37 0.25 ;
      LAYER M2 ;
      RECT 306.23 0.0 306.37 0.25 ;
      LAYER M3 ;
      RECT 306.23 0.0 306.37 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[42]
  PIN DB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 136.06 0.0 136.2 0.25 ;
      LAYER M2 ;
      RECT 136.06 0.0 136.2 0.25 ;
      LAYER M1 ;
      RECT 136.06 0.0 136.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[21]
  PIN DA[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 309.54 0.0 309.68 0.25 ;
      LAYER M2 ;
      RECT 309.54 0.0 309.68 0.25 ;
      LAYER M3 ;
      RECT 309.54 0.0 309.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[42]
  PIN DA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 132.75 0.0 132.89 0.25 ;
      LAYER M2 ;
      RECT 132.75 0.0 132.89 0.25 ;
      LAYER M1 ;
      RECT 132.75 0.0 132.89 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[21]
  PIN QA[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 310.325 0.0 310.465 0.25 ;
      LAYER M2 ;
      RECT 310.325 0.0 310.465 0.25 ;
      LAYER M3 ;
      RECT 310.325 0.0 310.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[42]
  PIN QA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 131.965 0.0 132.105 0.25 ;
      LAYER M2 ;
      RECT 131.965 0.0 132.105 0.25 ;
      LAYER M1 ;
      RECT 131.965 0.0 132.105 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[21]
  PIN TDA[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 310.705 0.0 310.845 0.25 ;
      LAYER M2 ;
      RECT 310.705 0.0 310.845 0.25 ;
      LAYER M3 ;
      RECT 310.705 0.0 310.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[42]
  PIN TDA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 131.585 0.0 131.725 0.25 ;
      LAYER M2 ;
      RECT 131.585 0.0 131.725 0.25 ;
      LAYER M1 ;
      RECT 131.585 0.0 131.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[21]
  PIN TDB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 311.27 0.0 311.41 0.25 ;
      LAYER M2 ;
      RECT 311.27 0.0 311.41 0.25 ;
      LAYER M3 ;
      RECT 311.27 0.0 311.41 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[43]
  PIN TDB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 131.02 0.0 131.16 0.25 ;
      LAYER M2 ;
      RECT 131.02 0.0 131.16 0.25 ;
      LAYER M1 ;
      RECT 131.02 0.0 131.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[20]
  PIN QB[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 311.655 0.0 311.795 0.25 ;
      LAYER M2 ;
      RECT 311.655 0.0 311.795 0.25 ;
      LAYER M3 ;
      RECT 311.655 0.0 311.795 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[43]
  PIN QB[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 130.635 0.0 130.775 0.25 ;
      LAYER M2 ;
      RECT 130.635 0.0 130.775 0.25 ;
      LAYER M1 ;
      RECT 130.635 0.0 130.775 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[20]
  PIN DB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 312.43 0.0 312.57 0.25 ;
      LAYER M2 ;
      RECT 312.43 0.0 312.57 0.25 ;
      LAYER M3 ;
      RECT 312.43 0.0 312.57 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[43]
  PIN DB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 129.86 0.0 130.0 0.25 ;
      LAYER M2 ;
      RECT 129.86 0.0 130.0 0.25 ;
      LAYER M1 ;
      RECT 129.86 0.0 130.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[20]
  PIN DA[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 315.74 0.0 315.88 0.25 ;
      LAYER M2 ;
      RECT 315.74 0.0 315.88 0.25 ;
      LAYER M3 ;
      RECT 315.74 0.0 315.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[43]
  PIN DA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 126.55 0.0 126.69 0.25 ;
      LAYER M2 ;
      RECT 126.55 0.0 126.69 0.25 ;
      LAYER M1 ;
      RECT 126.55 0.0 126.69 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[20]
  PIN QA[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 316.525 0.0 316.665 0.25 ;
      LAYER M2 ;
      RECT 316.525 0.0 316.665 0.25 ;
      LAYER M3 ;
      RECT 316.525 0.0 316.665 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[43]
  PIN QA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 125.765 0.0 125.905 0.25 ;
      LAYER M2 ;
      RECT 125.765 0.0 125.905 0.25 ;
      LAYER M1 ;
      RECT 125.765 0.0 125.905 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[20]
  PIN TDA[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 316.905 0.0 317.045 0.25 ;
      LAYER M2 ;
      RECT 316.905 0.0 317.045 0.25 ;
      LAYER M3 ;
      RECT 316.905 0.0 317.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[43]
  PIN TDA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 125.385 0.0 125.525 0.25 ;
      LAYER M2 ;
      RECT 125.385 0.0 125.525 0.25 ;
      LAYER M1 ;
      RECT 125.385 0.0 125.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[20]
  PIN TDB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 317.47 0.0 317.61 0.25 ;
      LAYER M2 ;
      RECT 317.47 0.0 317.61 0.25 ;
      LAYER M3 ;
      RECT 317.47 0.0 317.61 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[44]
  PIN TDB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 124.82 0.0 124.96 0.25 ;
      LAYER M2 ;
      RECT 124.82 0.0 124.96 0.25 ;
      LAYER M1 ;
      RECT 124.82 0.0 124.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[19]
  PIN QB[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 317.855 0.0 317.995 0.25 ;
      LAYER M2 ;
      RECT 317.855 0.0 317.995 0.25 ;
      LAYER M3 ;
      RECT 317.855 0.0 317.995 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[44]
  PIN QB[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 124.435 0.0 124.575 0.25 ;
      LAYER M2 ;
      RECT 124.435 0.0 124.575 0.25 ;
      LAYER M1 ;
      RECT 124.435 0.0 124.575 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[19]
  PIN DB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 318.63 0.0 318.77 0.25 ;
      LAYER M2 ;
      RECT 318.63 0.0 318.77 0.25 ;
      LAYER M3 ;
      RECT 318.63 0.0 318.77 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[44]
  PIN DB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 123.66 0.0 123.8 0.25 ;
      LAYER M2 ;
      RECT 123.66 0.0 123.8 0.25 ;
      LAYER M1 ;
      RECT 123.66 0.0 123.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[19]
  PIN DA[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 321.94 0.0 322.08 0.25 ;
      LAYER M2 ;
      RECT 321.94 0.0 322.08 0.25 ;
      LAYER M3 ;
      RECT 321.94 0.0 322.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[44]
  PIN DA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 120.35 0.0 120.49 0.25 ;
      LAYER M2 ;
      RECT 120.35 0.0 120.49 0.25 ;
      LAYER M1 ;
      RECT 120.35 0.0 120.49 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[19]
  PIN QA[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 322.725 0.0 322.865 0.25 ;
      LAYER M2 ;
      RECT 322.725 0.0 322.865 0.25 ;
      LAYER M3 ;
      RECT 322.725 0.0 322.865 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[44]
  PIN QA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 119.565 0.0 119.705 0.25 ;
      LAYER M2 ;
      RECT 119.565 0.0 119.705 0.25 ;
      LAYER M1 ;
      RECT 119.565 0.0 119.705 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[19]
  PIN TDA[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 323.105 0.0 323.245 0.25 ;
      LAYER M2 ;
      RECT 323.105 0.0 323.245 0.25 ;
      LAYER M3 ;
      RECT 323.105 0.0 323.245 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[44]
  PIN TDA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 119.185 0.0 119.325 0.25 ;
      LAYER M2 ;
      RECT 119.185 0.0 119.325 0.25 ;
      LAYER M1 ;
      RECT 119.185 0.0 119.325 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[19]
  PIN TDB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 323.67 0.0 323.81 0.25 ;
      LAYER M2 ;
      RECT 323.67 0.0 323.81 0.25 ;
      LAYER M3 ;
      RECT 323.67 0.0 323.81 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[45]
  PIN TDB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.62 0.0 118.76 0.25 ;
      LAYER M2 ;
      RECT 118.62 0.0 118.76 0.25 ;
      LAYER M1 ;
      RECT 118.62 0.0 118.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[18]
  PIN QB[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 324.055 0.0 324.195 0.25 ;
      LAYER M2 ;
      RECT 324.055 0.0 324.195 0.25 ;
      LAYER M3 ;
      RECT 324.055 0.0 324.195 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[45]
  PIN QB[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 118.235 0.0 118.375 0.25 ;
      LAYER M2 ;
      RECT 118.235 0.0 118.375 0.25 ;
      LAYER M1 ;
      RECT 118.235 0.0 118.375 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[18]
  PIN DB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 324.83 0.0 324.97 0.25 ;
      LAYER M2 ;
      RECT 324.83 0.0 324.97 0.25 ;
      LAYER M3 ;
      RECT 324.83 0.0 324.97 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[45]
  PIN DB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 117.46 0.0 117.6 0.25 ;
      LAYER M2 ;
      RECT 117.46 0.0 117.6 0.25 ;
      LAYER M1 ;
      RECT 117.46 0.0 117.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[18]
  PIN DA[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 328.14 0.0 328.28 0.25 ;
      LAYER M2 ;
      RECT 328.14 0.0 328.28 0.25 ;
      LAYER M3 ;
      RECT 328.14 0.0 328.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[45]
  PIN DA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 114.15 0.0 114.29 0.25 ;
      LAYER M2 ;
      RECT 114.15 0.0 114.29 0.25 ;
      LAYER M1 ;
      RECT 114.15 0.0 114.29 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[18]
  PIN QA[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 328.925 0.0 329.065 0.25 ;
      LAYER M2 ;
      RECT 328.925 0.0 329.065 0.25 ;
      LAYER M3 ;
      RECT 328.925 0.0 329.065 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[45]
  PIN QA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 113.365 0.0 113.505 0.25 ;
      LAYER M2 ;
      RECT 113.365 0.0 113.505 0.25 ;
      LAYER M1 ;
      RECT 113.365 0.0 113.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[18]
  PIN TDA[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 329.305 0.0 329.445 0.25 ;
      LAYER M2 ;
      RECT 329.305 0.0 329.445 0.25 ;
      LAYER M3 ;
      RECT 329.305 0.0 329.445 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[45]
  PIN TDA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 112.985 0.0 113.125 0.25 ;
      LAYER M2 ;
      RECT 112.985 0.0 113.125 0.25 ;
      LAYER M1 ;
      RECT 112.985 0.0 113.125 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[18]
  PIN TDB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 329.87 0.0 330.01 0.25 ;
      LAYER M2 ;
      RECT 329.87 0.0 330.01 0.25 ;
      LAYER M3 ;
      RECT 329.87 0.0 330.01 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[46]
  PIN TDB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 112.42 0.0 112.56 0.25 ;
      LAYER M2 ;
      RECT 112.42 0.0 112.56 0.25 ;
      LAYER M1 ;
      RECT 112.42 0.0 112.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[17]
  PIN QB[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 330.255 0.0 330.395 0.25 ;
      LAYER M2 ;
      RECT 330.255 0.0 330.395 0.25 ;
      LAYER M3 ;
      RECT 330.255 0.0 330.395 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[46]
  PIN QB[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 112.035 0.0 112.175 0.25 ;
      LAYER M2 ;
      RECT 112.035 0.0 112.175 0.25 ;
      LAYER M1 ;
      RECT 112.035 0.0 112.175 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[17]
  PIN DB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 331.03 0.0 331.17 0.25 ;
      LAYER M2 ;
      RECT 331.03 0.0 331.17 0.25 ;
      LAYER M3 ;
      RECT 331.03 0.0 331.17 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[46]
  PIN DB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 111.26 0.0 111.4 0.25 ;
      LAYER M2 ;
      RECT 111.26 0.0 111.4 0.25 ;
      LAYER M1 ;
      RECT 111.26 0.0 111.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[17]
  PIN DA[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 334.34 0.0 334.48 0.25 ;
      LAYER M2 ;
      RECT 334.34 0.0 334.48 0.25 ;
      LAYER M3 ;
      RECT 334.34 0.0 334.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[46]
  PIN DA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 107.95 0.0 108.09 0.25 ;
      LAYER M2 ;
      RECT 107.95 0.0 108.09 0.25 ;
      LAYER M1 ;
      RECT 107.95 0.0 108.09 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[17]
  PIN QA[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 335.125 0.0 335.265 0.25 ;
      LAYER M2 ;
      RECT 335.125 0.0 335.265 0.25 ;
      LAYER M3 ;
      RECT 335.125 0.0 335.265 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[46]
  PIN QA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 107.165 0.0 107.305 0.25 ;
      LAYER M2 ;
      RECT 107.165 0.0 107.305 0.25 ;
      LAYER M1 ;
      RECT 107.165 0.0 107.305 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[17]
  PIN TDA[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 335.505 0.0 335.645 0.25 ;
      LAYER M2 ;
      RECT 335.505 0.0 335.645 0.25 ;
      LAYER M3 ;
      RECT 335.505 0.0 335.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[46]
  PIN TDA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 106.785 0.0 106.925 0.25 ;
      LAYER M2 ;
      RECT 106.785 0.0 106.925 0.25 ;
      LAYER M1 ;
      RECT 106.785 0.0 106.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[17]
  PIN TDB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 336.07 0.0 336.21 0.25 ;
      LAYER M2 ;
      RECT 336.07 0.0 336.21 0.25 ;
      LAYER M3 ;
      RECT 336.07 0.0 336.21 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[47]
  PIN TDB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 106.22 0.0 106.36 0.25 ;
      LAYER M2 ;
      RECT 106.22 0.0 106.36 0.25 ;
      LAYER M1 ;
      RECT 106.22 0.0 106.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[16]
  PIN QB[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 336.455 0.0 336.595 0.25 ;
      LAYER M2 ;
      RECT 336.455 0.0 336.595 0.25 ;
      LAYER M3 ;
      RECT 336.455 0.0 336.595 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[47]
  PIN QB[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 105.835 0.0 105.975 0.25 ;
      LAYER M2 ;
      RECT 105.835 0.0 105.975 0.25 ;
      LAYER M1 ;
      RECT 105.835 0.0 105.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[16]
  PIN DB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 337.23 0.0 337.37 0.25 ;
      LAYER M2 ;
      RECT 337.23 0.0 337.37 0.25 ;
      LAYER M3 ;
      RECT 337.23 0.0 337.37 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[47]
  PIN DB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 105.06 0.0 105.2 0.25 ;
      LAYER M2 ;
      RECT 105.06 0.0 105.2 0.25 ;
      LAYER M1 ;
      RECT 105.06 0.0 105.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[16]
  PIN DA[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 340.54 0.0 340.68 0.25 ;
      LAYER M2 ;
      RECT 340.54 0.0 340.68 0.25 ;
      LAYER M3 ;
      RECT 340.54 0.0 340.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[47]
  PIN DA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 101.75 0.0 101.89 0.25 ;
      LAYER M2 ;
      RECT 101.75 0.0 101.89 0.25 ;
      LAYER M1 ;
      RECT 101.75 0.0 101.89 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[16]
  PIN QA[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 341.325 0.0 341.465 0.25 ;
      LAYER M2 ;
      RECT 341.325 0.0 341.465 0.25 ;
      LAYER M3 ;
      RECT 341.325 0.0 341.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[47]
  PIN QA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 100.965 0.0 101.105 0.25 ;
      LAYER M2 ;
      RECT 100.965 0.0 101.105 0.25 ;
      LAYER M1 ;
      RECT 100.965 0.0 101.105 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[16]
  PIN TDA[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 341.705 0.0 341.845 0.25 ;
      LAYER M2 ;
      RECT 341.705 0.0 341.845 0.25 ;
      LAYER M3 ;
      RECT 341.705 0.0 341.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[47]
  PIN TDA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 100.585 0.0 100.725 0.25 ;
      LAYER M2 ;
      RECT 100.585 0.0 100.725 0.25 ;
      LAYER M1 ;
      RECT 100.585 0.0 100.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[16]
  PIN TDB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 342.27 0.0 342.41 0.25 ;
      LAYER M2 ;
      RECT 342.27 0.0 342.41 0.25 ;
      LAYER M3 ;
      RECT 342.27 0.0 342.41 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[48]
  PIN TDB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 100.02 0.0 100.16 0.25 ;
      LAYER M2 ;
      RECT 100.02 0.0 100.16 0.25 ;
      LAYER M1 ;
      RECT 100.02 0.0 100.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[15]
  PIN QB[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 342.655 0.0 342.795 0.25 ;
      LAYER M2 ;
      RECT 342.655 0.0 342.795 0.25 ;
      LAYER M3 ;
      RECT 342.655 0.0 342.795 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[48]
  PIN QB[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 99.635 0.0 99.775 0.25 ;
      LAYER M2 ;
      RECT 99.635 0.0 99.775 0.25 ;
      LAYER M1 ;
      RECT 99.635 0.0 99.775 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[15]
  PIN DB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 343.43 0.0 343.57 0.25 ;
      LAYER M2 ;
      RECT 343.43 0.0 343.57 0.25 ;
      LAYER M3 ;
      RECT 343.43 0.0 343.57 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[48]
  PIN DB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 98.86 0.0 99.0 0.25 ;
      LAYER M2 ;
      RECT 98.86 0.0 99.0 0.25 ;
      LAYER M1 ;
      RECT 98.86 0.0 99.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[15]
  PIN DA[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 346.74 0.0 346.88 0.25 ;
      LAYER M2 ;
      RECT 346.74 0.0 346.88 0.25 ;
      LAYER M3 ;
      RECT 346.74 0.0 346.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[48]
  PIN DA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 95.55 0.0 95.69 0.25 ;
      LAYER M2 ;
      RECT 95.55 0.0 95.69 0.25 ;
      LAYER M1 ;
      RECT 95.55 0.0 95.69 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[15]
  PIN QA[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 347.525 0.0 347.665 0.25 ;
      LAYER M2 ;
      RECT 347.525 0.0 347.665 0.25 ;
      LAYER M3 ;
      RECT 347.525 0.0 347.665 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[48]
  PIN QA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 94.765 0.0 94.905 0.25 ;
      LAYER M2 ;
      RECT 94.765 0.0 94.905 0.25 ;
      LAYER M1 ;
      RECT 94.765 0.0 94.905 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[15]
  PIN TDA[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 347.905 0.0 348.045 0.25 ;
      LAYER M2 ;
      RECT 347.905 0.0 348.045 0.25 ;
      LAYER M3 ;
      RECT 347.905 0.0 348.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[48]
  PIN TDA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 94.385 0.0 94.525 0.25 ;
      LAYER M2 ;
      RECT 94.385 0.0 94.525 0.25 ;
      LAYER M1 ;
      RECT 94.385 0.0 94.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[15]
  PIN TDB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 348.47 0.0 348.61 0.25 ;
      LAYER M2 ;
      RECT 348.47 0.0 348.61 0.25 ;
      LAYER M3 ;
      RECT 348.47 0.0 348.61 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[49]
  PIN TDB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 93.82 0.0 93.96 0.25 ;
      LAYER M2 ;
      RECT 93.82 0.0 93.96 0.25 ;
      LAYER M1 ;
      RECT 93.82 0.0 93.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[14]
  PIN QB[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 348.855 0.0 348.995 0.25 ;
      LAYER M2 ;
      RECT 348.855 0.0 348.995 0.25 ;
      LAYER M3 ;
      RECT 348.855 0.0 348.995 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[49]
  PIN QB[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 93.435 0.0 93.575 0.25 ;
      LAYER M2 ;
      RECT 93.435 0.0 93.575 0.25 ;
      LAYER M1 ;
      RECT 93.435 0.0 93.575 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[14]
  PIN DB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 349.63 0.0 349.77 0.25 ;
      LAYER M2 ;
      RECT 349.63 0.0 349.77 0.25 ;
      LAYER M3 ;
      RECT 349.63 0.0 349.77 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[49]
  PIN DB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 92.66 0.0 92.8 0.25 ;
      LAYER M2 ;
      RECT 92.66 0.0 92.8 0.25 ;
      LAYER M1 ;
      RECT 92.66 0.0 92.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[14]
  PIN DA[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 352.94 0.0 353.08 0.25 ;
      LAYER M2 ;
      RECT 352.94 0.0 353.08 0.25 ;
      LAYER M3 ;
      RECT 352.94 0.0 353.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[49]
  PIN DA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 89.35 0.0 89.49 0.25 ;
      LAYER M2 ;
      RECT 89.35 0.0 89.49 0.25 ;
      LAYER M1 ;
      RECT 89.35 0.0 89.49 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[14]
  PIN QA[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 353.725 0.0 353.865 0.25 ;
      LAYER M2 ;
      RECT 353.725 0.0 353.865 0.25 ;
      LAYER M3 ;
      RECT 353.725 0.0 353.865 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[49]
  PIN QA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.565 0.0 88.705 0.25 ;
      LAYER M2 ;
      RECT 88.565 0.0 88.705 0.25 ;
      LAYER M1 ;
      RECT 88.565 0.0 88.705 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[14]
  PIN TDA[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 354.105 0.0 354.245 0.25 ;
      LAYER M2 ;
      RECT 354.105 0.0 354.245 0.25 ;
      LAYER M3 ;
      RECT 354.105 0.0 354.245 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[49]
  PIN TDA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 88.185 0.0 88.325 0.25 ;
      LAYER M2 ;
      RECT 88.185 0.0 88.325 0.25 ;
      LAYER M1 ;
      RECT 88.185 0.0 88.325 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[14]
  PIN TDB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 354.67 0.0 354.81 0.25 ;
      LAYER M2 ;
      RECT 354.67 0.0 354.81 0.25 ;
      LAYER M3 ;
      RECT 354.67 0.0 354.81 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[50]
  PIN TDB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 87.62 0.0 87.76 0.25 ;
      LAYER M2 ;
      RECT 87.62 0.0 87.76 0.25 ;
      LAYER M1 ;
      RECT 87.62 0.0 87.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[13]
  PIN QB[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 355.055 0.0 355.195 0.25 ;
      LAYER M2 ;
      RECT 355.055 0.0 355.195 0.25 ;
      LAYER M3 ;
      RECT 355.055 0.0 355.195 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[50]
  PIN QB[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 87.235 0.0 87.375 0.25 ;
      LAYER M2 ;
      RECT 87.235 0.0 87.375 0.25 ;
      LAYER M1 ;
      RECT 87.235 0.0 87.375 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[13]
  PIN DB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 355.83 0.0 355.97 0.25 ;
      LAYER M2 ;
      RECT 355.83 0.0 355.97 0.25 ;
      LAYER M3 ;
      RECT 355.83 0.0 355.97 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[50]
  PIN DB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 86.46 0.0 86.6 0.25 ;
      LAYER M2 ;
      RECT 86.46 0.0 86.6 0.25 ;
      LAYER M1 ;
      RECT 86.46 0.0 86.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[13]
  PIN DA[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 359.14 0.0 359.28 0.25 ;
      LAYER M2 ;
      RECT 359.14 0.0 359.28 0.25 ;
      LAYER M3 ;
      RECT 359.14 0.0 359.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[50]
  PIN DA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 83.15 0.0 83.29 0.25 ;
      LAYER M2 ;
      RECT 83.15 0.0 83.29 0.25 ;
      LAYER M1 ;
      RECT 83.15 0.0 83.29 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[13]
  PIN QA[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 359.925 0.0 360.065 0.25 ;
      LAYER M2 ;
      RECT 359.925 0.0 360.065 0.25 ;
      LAYER M3 ;
      RECT 359.925 0.0 360.065 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[50]
  PIN QA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 82.365 0.0 82.505 0.25 ;
      LAYER M2 ;
      RECT 82.365 0.0 82.505 0.25 ;
      LAYER M1 ;
      RECT 82.365 0.0 82.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[13]
  PIN TDA[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 360.305 0.0 360.445 0.25 ;
      LAYER M2 ;
      RECT 360.305 0.0 360.445 0.25 ;
      LAYER M3 ;
      RECT 360.305 0.0 360.445 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[50]
  PIN TDA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 81.985 0.0 82.125 0.25 ;
      LAYER M2 ;
      RECT 81.985 0.0 82.125 0.25 ;
      LAYER M1 ;
      RECT 81.985 0.0 82.125 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[13]
  PIN TDB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 360.87 0.0 361.01 0.25 ;
      LAYER M2 ;
      RECT 360.87 0.0 361.01 0.25 ;
      LAYER M3 ;
      RECT 360.87 0.0 361.01 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[51]
  PIN TDB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 81.42 0.0 81.56 0.25 ;
      LAYER M2 ;
      RECT 81.42 0.0 81.56 0.25 ;
      LAYER M1 ;
      RECT 81.42 0.0 81.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[12]
  PIN QB[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 361.255 0.0 361.395 0.25 ;
      LAYER M2 ;
      RECT 361.255 0.0 361.395 0.25 ;
      LAYER M3 ;
      RECT 361.255 0.0 361.395 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[51]
  PIN QB[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 81.035 0.0 81.175 0.25 ;
      LAYER M2 ;
      RECT 81.035 0.0 81.175 0.25 ;
      LAYER M1 ;
      RECT 81.035 0.0 81.175 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[12]
  PIN DB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 362.03 0.0 362.17 0.25 ;
      LAYER M2 ;
      RECT 362.03 0.0 362.17 0.25 ;
      LAYER M3 ;
      RECT 362.03 0.0 362.17 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[51]
  PIN DB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 80.26 0.0 80.4 0.25 ;
      LAYER M2 ;
      RECT 80.26 0.0 80.4 0.25 ;
      LAYER M1 ;
      RECT 80.26 0.0 80.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[12]
  PIN DA[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 365.34 0.0 365.48 0.25 ;
      LAYER M2 ;
      RECT 365.34 0.0 365.48 0.25 ;
      LAYER M3 ;
      RECT 365.34 0.0 365.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[51]
  PIN DA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 76.95 0.0 77.09 0.25 ;
      LAYER M2 ;
      RECT 76.95 0.0 77.09 0.25 ;
      LAYER M1 ;
      RECT 76.95 0.0 77.09 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[12]
  PIN QA[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 366.125 0.0 366.265 0.25 ;
      LAYER M2 ;
      RECT 366.125 0.0 366.265 0.25 ;
      LAYER M3 ;
      RECT 366.125 0.0 366.265 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[51]
  PIN QA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 76.165 0.0 76.305 0.25 ;
      LAYER M2 ;
      RECT 76.165 0.0 76.305 0.25 ;
      LAYER M1 ;
      RECT 76.165 0.0 76.305 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[12]
  PIN TDA[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 366.505 0.0 366.645 0.25 ;
      LAYER M2 ;
      RECT 366.505 0.0 366.645 0.25 ;
      LAYER M3 ;
      RECT 366.505 0.0 366.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[51]
  PIN TDA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 75.785 0.0 75.925 0.25 ;
      LAYER M2 ;
      RECT 75.785 0.0 75.925 0.25 ;
      LAYER M1 ;
      RECT 75.785 0.0 75.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[12]
  PIN TDB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 367.07 0.0 367.21 0.25 ;
      LAYER M2 ;
      RECT 367.07 0.0 367.21 0.25 ;
      LAYER M3 ;
      RECT 367.07 0.0 367.21 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[52]
  PIN TDB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 75.22 0.0 75.36 0.25 ;
      LAYER M2 ;
      RECT 75.22 0.0 75.36 0.25 ;
      LAYER M1 ;
      RECT 75.22 0.0 75.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[11]
  PIN QB[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 367.455 0.0 367.595 0.25 ;
      LAYER M2 ;
      RECT 367.455 0.0 367.595 0.25 ;
      LAYER M3 ;
      RECT 367.455 0.0 367.595 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[52]
  PIN QB[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 74.835 0.0 74.975 0.25 ;
      LAYER M2 ;
      RECT 74.835 0.0 74.975 0.25 ;
      LAYER M1 ;
      RECT 74.835 0.0 74.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[11]
  PIN DB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 368.23 0.0 368.37 0.25 ;
      LAYER M2 ;
      RECT 368.23 0.0 368.37 0.25 ;
      LAYER M3 ;
      RECT 368.23 0.0 368.37 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[52]
  PIN DB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 74.06 0.0 74.2 0.25 ;
      LAYER M2 ;
      RECT 74.06 0.0 74.2 0.25 ;
      LAYER M1 ;
      RECT 74.06 0.0 74.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[11]
  PIN DA[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 371.54 0.0 371.68 0.25 ;
      LAYER M2 ;
      RECT 371.54 0.0 371.68 0.25 ;
      LAYER M3 ;
      RECT 371.54 0.0 371.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[52]
  PIN DA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 70.75 0.0 70.89 0.25 ;
      LAYER M2 ;
      RECT 70.75 0.0 70.89 0.25 ;
      LAYER M1 ;
      RECT 70.75 0.0 70.89 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[11]
  PIN QA[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 372.325 0.0 372.465 0.25 ;
      LAYER M2 ;
      RECT 372.325 0.0 372.465 0.25 ;
      LAYER M3 ;
      RECT 372.325 0.0 372.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[52]
  PIN QA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.965 0.0 70.105 0.25 ;
      LAYER M2 ;
      RECT 69.965 0.0 70.105 0.25 ;
      LAYER M1 ;
      RECT 69.965 0.0 70.105 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[11]
  PIN TDA[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 372.705 0.0 372.845 0.25 ;
      LAYER M2 ;
      RECT 372.705 0.0 372.845 0.25 ;
      LAYER M3 ;
      RECT 372.705 0.0 372.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[52]
  PIN TDA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.585 0.0 69.725 0.25 ;
      LAYER M2 ;
      RECT 69.585 0.0 69.725 0.25 ;
      LAYER M1 ;
      RECT 69.585 0.0 69.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[11]
  PIN TDB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 373.27 0.0 373.41 0.25 ;
      LAYER M2 ;
      RECT 373.27 0.0 373.41 0.25 ;
      LAYER M3 ;
      RECT 373.27 0.0 373.41 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[53]
  PIN TDB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 69.02 0.0 69.16 0.25 ;
      LAYER M2 ;
      RECT 69.02 0.0 69.16 0.25 ;
      LAYER M1 ;
      RECT 69.02 0.0 69.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[10]
  PIN QB[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 373.655 0.0 373.795 0.25 ;
      LAYER M2 ;
      RECT 373.655 0.0 373.795 0.25 ;
      LAYER M3 ;
      RECT 373.655 0.0 373.795 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[53]
  PIN QB[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 68.635 0.0 68.775 0.25 ;
      LAYER M2 ;
      RECT 68.635 0.0 68.775 0.25 ;
      LAYER M1 ;
      RECT 68.635 0.0 68.775 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[10]
  PIN DB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 374.43 0.0 374.57 0.25 ;
      LAYER M2 ;
      RECT 374.43 0.0 374.57 0.25 ;
      LAYER M3 ;
      RECT 374.43 0.0 374.57 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[53]
  PIN DB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 67.86 0.0 68.0 0.25 ;
      LAYER M2 ;
      RECT 67.86 0.0 68.0 0.25 ;
      LAYER M1 ;
      RECT 67.86 0.0 68.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[10]
  PIN DA[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 377.74 0.0 377.88 0.25 ;
      LAYER M2 ;
      RECT 377.74 0.0 377.88 0.25 ;
      LAYER M3 ;
      RECT 377.74 0.0 377.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[53]
  PIN DA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 64.55 0.0 64.69 0.25 ;
      LAYER M2 ;
      RECT 64.55 0.0 64.69 0.25 ;
      LAYER M1 ;
      RECT 64.55 0.0 64.69 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[10]
  PIN QA[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 378.525 0.0 378.665 0.25 ;
      LAYER M2 ;
      RECT 378.525 0.0 378.665 0.25 ;
      LAYER M3 ;
      RECT 378.525 0.0 378.665 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[53]
  PIN QA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 63.765 0.0 63.905 0.25 ;
      LAYER M2 ;
      RECT 63.765 0.0 63.905 0.25 ;
      LAYER M1 ;
      RECT 63.765 0.0 63.905 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[10]
  PIN TDA[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 378.905 0.0 379.045 0.25 ;
      LAYER M2 ;
      RECT 378.905 0.0 379.045 0.25 ;
      LAYER M3 ;
      RECT 378.905 0.0 379.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[53]
  PIN TDA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 63.385 0.0 63.525 0.25 ;
      LAYER M2 ;
      RECT 63.385 0.0 63.525 0.25 ;
      LAYER M1 ;
      RECT 63.385 0.0 63.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[10]
  PIN TDB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 379.47 0.0 379.61 0.25 ;
      LAYER M2 ;
      RECT 379.47 0.0 379.61 0.25 ;
      LAYER M3 ;
      RECT 379.47 0.0 379.61 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[54]
  PIN TDB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 62.82 0.0 62.96 0.25 ;
      LAYER M2 ;
      RECT 62.82 0.0 62.96 0.25 ;
      LAYER M1 ;
      RECT 62.82 0.0 62.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[9]
  PIN QB[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 379.855 0.0 379.995 0.25 ;
      LAYER M2 ;
      RECT 379.855 0.0 379.995 0.25 ;
      LAYER M3 ;
      RECT 379.855 0.0 379.995 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[54]
  PIN QB[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 62.435 0.0 62.575 0.25 ;
      LAYER M2 ;
      RECT 62.435 0.0 62.575 0.25 ;
      LAYER M1 ;
      RECT 62.435 0.0 62.575 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[9]
  PIN DB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 380.63 0.0 380.77 0.25 ;
      LAYER M2 ;
      RECT 380.63 0.0 380.77 0.25 ;
      LAYER M3 ;
      RECT 380.63 0.0 380.77 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[54]
  PIN DB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 61.66 0.0 61.8 0.25 ;
      LAYER M2 ;
      RECT 61.66 0.0 61.8 0.25 ;
      LAYER M1 ;
      RECT 61.66 0.0 61.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[9]
  PIN DA[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 383.94 0.0 384.08 0.25 ;
      LAYER M2 ;
      RECT 383.94 0.0 384.08 0.25 ;
      LAYER M3 ;
      RECT 383.94 0.0 384.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[54]
  PIN DA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 58.35 0.0 58.49 0.25 ;
      LAYER M2 ;
      RECT 58.35 0.0 58.49 0.25 ;
      LAYER M1 ;
      RECT 58.35 0.0 58.49 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[9]
  PIN QA[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 384.725 0.0 384.865 0.25 ;
      LAYER M2 ;
      RECT 384.725 0.0 384.865 0.25 ;
      LAYER M3 ;
      RECT 384.725 0.0 384.865 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[54]
  PIN QA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 57.565 0.0 57.705 0.25 ;
      LAYER M2 ;
      RECT 57.565 0.0 57.705 0.25 ;
      LAYER M1 ;
      RECT 57.565 0.0 57.705 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[9]
  PIN TDA[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 385.105 0.0 385.245 0.25 ;
      LAYER M2 ;
      RECT 385.105 0.0 385.245 0.25 ;
      LAYER M3 ;
      RECT 385.105 0.0 385.245 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[54]
  PIN TDA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 57.185 0.0 57.325 0.25 ;
      LAYER M2 ;
      RECT 57.185 0.0 57.325 0.25 ;
      LAYER M1 ;
      RECT 57.185 0.0 57.325 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[9]
  PIN TDB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 385.67 0.0 385.81 0.25 ;
      LAYER M2 ;
      RECT 385.67 0.0 385.81 0.25 ;
      LAYER M3 ;
      RECT 385.67 0.0 385.81 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[55]
  PIN TDB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 56.62 0.0 56.76 0.25 ;
      LAYER M2 ;
      RECT 56.62 0.0 56.76 0.25 ;
      LAYER M1 ;
      RECT 56.62 0.0 56.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[8]
  PIN QB[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 386.055 0.0 386.195 0.25 ;
      LAYER M2 ;
      RECT 386.055 0.0 386.195 0.25 ;
      LAYER M3 ;
      RECT 386.055 0.0 386.195 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[55]
  PIN QB[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 56.235 0.0 56.375 0.25 ;
      LAYER M2 ;
      RECT 56.235 0.0 56.375 0.25 ;
      LAYER M1 ;
      RECT 56.235 0.0 56.375 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[8]
  PIN DB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 386.83 0.0 386.97 0.25 ;
      LAYER M2 ;
      RECT 386.83 0.0 386.97 0.25 ;
      LAYER M3 ;
      RECT 386.83 0.0 386.97 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[55]
  PIN DB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 55.46 0.0 55.6 0.25 ;
      LAYER M2 ;
      RECT 55.46 0.0 55.6 0.25 ;
      LAYER M1 ;
      RECT 55.46 0.0 55.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[8]
  PIN DA[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 390.14 0.0 390.28 0.25 ;
      LAYER M2 ;
      RECT 390.14 0.0 390.28 0.25 ;
      LAYER M3 ;
      RECT 390.14 0.0 390.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[55]
  PIN DA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 52.15 0.0 52.29 0.25 ;
      LAYER M2 ;
      RECT 52.15 0.0 52.29 0.25 ;
      LAYER M1 ;
      RECT 52.15 0.0 52.29 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[8]
  PIN QA[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 390.925 0.0 391.065 0.25 ;
      LAYER M2 ;
      RECT 390.925 0.0 391.065 0.25 ;
      LAYER M3 ;
      RECT 390.925 0.0 391.065 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[55]
  PIN QA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 51.365 0.0 51.505 0.25 ;
      LAYER M2 ;
      RECT 51.365 0.0 51.505 0.25 ;
      LAYER M1 ;
      RECT 51.365 0.0 51.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[8]
  PIN TDA[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 391.305 0.0 391.445 0.25 ;
      LAYER M2 ;
      RECT 391.305 0.0 391.445 0.25 ;
      LAYER M3 ;
      RECT 391.305 0.0 391.445 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[55]
  PIN TDA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 50.985 0.0 51.125 0.25 ;
      LAYER M2 ;
      RECT 50.985 0.0 51.125 0.25 ;
      LAYER M1 ;
      RECT 50.985 0.0 51.125 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[8]
  PIN TDB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 391.87 0.0 392.01 0.25 ;
      LAYER M2 ;
      RECT 391.87 0.0 392.01 0.25 ;
      LAYER M3 ;
      RECT 391.87 0.0 392.01 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[56]
  PIN TDB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 50.42 0.0 50.56 0.25 ;
      LAYER M2 ;
      RECT 50.42 0.0 50.56 0.25 ;
      LAYER M1 ;
      RECT 50.42 0.0 50.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[7]
  PIN QB[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 392.255 0.0 392.395 0.25 ;
      LAYER M2 ;
      RECT 392.255 0.0 392.395 0.25 ;
      LAYER M3 ;
      RECT 392.255 0.0 392.395 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[56]
  PIN QB[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 50.035 0.0 50.175 0.25 ;
      LAYER M2 ;
      RECT 50.035 0.0 50.175 0.25 ;
      LAYER M1 ;
      RECT 50.035 0.0 50.175 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[7]
  PIN DB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 393.03 0.0 393.17 0.25 ;
      LAYER M2 ;
      RECT 393.03 0.0 393.17 0.25 ;
      LAYER M3 ;
      RECT 393.03 0.0 393.17 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[56]
  PIN DB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.26 0.0 49.4 0.25 ;
      LAYER M2 ;
      RECT 49.26 0.0 49.4 0.25 ;
      LAYER M1 ;
      RECT 49.26 0.0 49.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[7]
  PIN DA[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 396.34 0.0 396.48 0.25 ;
      LAYER M2 ;
      RECT 396.34 0.0 396.48 0.25 ;
      LAYER M3 ;
      RECT 396.34 0.0 396.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[56]
  PIN DA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.95 0.0 46.09 0.25 ;
      LAYER M2 ;
      RECT 45.95 0.0 46.09 0.25 ;
      LAYER M1 ;
      RECT 45.95 0.0 46.09 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[7]
  PIN QA[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 397.125 0.0 397.265 0.25 ;
      LAYER M2 ;
      RECT 397.125 0.0 397.265 0.25 ;
      LAYER M3 ;
      RECT 397.125 0.0 397.265 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[56]
  PIN QA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.165 0.0 45.305 0.25 ;
      LAYER M2 ;
      RECT 45.165 0.0 45.305 0.25 ;
      LAYER M1 ;
      RECT 45.165 0.0 45.305 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[7]
  PIN TDA[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 397.505 0.0 397.645 0.25 ;
      LAYER M2 ;
      RECT 397.505 0.0 397.645 0.25 ;
      LAYER M3 ;
      RECT 397.505 0.0 397.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[56]
  PIN TDA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 44.785 0.0 44.925 0.25 ;
      LAYER M2 ;
      RECT 44.785 0.0 44.925 0.25 ;
      LAYER M1 ;
      RECT 44.785 0.0 44.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[7]
  PIN TDB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 398.07 0.0 398.21 0.25 ;
      LAYER M2 ;
      RECT 398.07 0.0 398.21 0.25 ;
      LAYER M3 ;
      RECT 398.07 0.0 398.21 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[57]
  PIN TDB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 44.22 0.0 44.36 0.25 ;
      LAYER M2 ;
      RECT 44.22 0.0 44.36 0.25 ;
      LAYER M1 ;
      RECT 44.22 0.0 44.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[6]
  PIN QB[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 398.455 0.0 398.595 0.25 ;
      LAYER M2 ;
      RECT 398.455 0.0 398.595 0.25 ;
      LAYER M3 ;
      RECT 398.455 0.0 398.595 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[57]
  PIN QB[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.835 0.0 43.975 0.25 ;
      LAYER M2 ;
      RECT 43.835 0.0 43.975 0.25 ;
      LAYER M1 ;
      RECT 43.835 0.0 43.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[6]
  PIN DB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 399.23 0.0 399.37 0.25 ;
      LAYER M2 ;
      RECT 399.23 0.0 399.37 0.25 ;
      LAYER M3 ;
      RECT 399.23 0.0 399.37 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[57]
  PIN DB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.06 0.0 43.2 0.25 ;
      LAYER M2 ;
      RECT 43.06 0.0 43.2 0.25 ;
      LAYER M1 ;
      RECT 43.06 0.0 43.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[6]
  PIN DA[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 402.54 0.0 402.68 0.25 ;
      LAYER M2 ;
      RECT 402.54 0.0 402.68 0.25 ;
      LAYER M3 ;
      RECT 402.54 0.0 402.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[57]
  PIN DA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.75 0.0 39.89 0.25 ;
      LAYER M2 ;
      RECT 39.75 0.0 39.89 0.25 ;
      LAYER M1 ;
      RECT 39.75 0.0 39.89 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[6]
  PIN QA[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 403.325 0.0 403.465 0.25 ;
      LAYER M2 ;
      RECT 403.325 0.0 403.465 0.25 ;
      LAYER M3 ;
      RECT 403.325 0.0 403.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[57]
  PIN QA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.965 0.0 39.105 0.25 ;
      LAYER M2 ;
      RECT 38.965 0.0 39.105 0.25 ;
      LAYER M1 ;
      RECT 38.965 0.0 39.105 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[6]
  PIN TDA[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 403.705 0.0 403.845 0.25 ;
      LAYER M2 ;
      RECT 403.705 0.0 403.845 0.25 ;
      LAYER M3 ;
      RECT 403.705 0.0 403.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[57]
  PIN TDA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.585 0.0 38.725 0.25 ;
      LAYER M2 ;
      RECT 38.585 0.0 38.725 0.25 ;
      LAYER M1 ;
      RECT 38.585 0.0 38.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[6]
  PIN TDB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 404.27 0.0 404.41 0.25 ;
      LAYER M2 ;
      RECT 404.27 0.0 404.41 0.25 ;
      LAYER M3 ;
      RECT 404.27 0.0 404.41 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[58]
  PIN TDB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.02 0.0 38.16 0.25 ;
      LAYER M2 ;
      RECT 38.02 0.0 38.16 0.25 ;
      LAYER M1 ;
      RECT 38.02 0.0 38.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[5]
  PIN QB[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 404.655 0.0 404.795 0.25 ;
      LAYER M2 ;
      RECT 404.655 0.0 404.795 0.25 ;
      LAYER M3 ;
      RECT 404.655 0.0 404.795 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[58]
  PIN QB[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 37.635 0.0 37.775 0.25 ;
      LAYER M2 ;
      RECT 37.635 0.0 37.775 0.25 ;
      LAYER M1 ;
      RECT 37.635 0.0 37.775 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[5]
  PIN DB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 405.43 0.0 405.57 0.25 ;
      LAYER M2 ;
      RECT 405.43 0.0 405.57 0.25 ;
      LAYER M3 ;
      RECT 405.43 0.0 405.57 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[58]
  PIN DB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 36.86 0.0 37.0 0.25 ;
      LAYER M2 ;
      RECT 36.86 0.0 37.0 0.25 ;
      LAYER M1 ;
      RECT 36.86 0.0 37.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[5]
  PIN DA[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 408.74 0.0 408.88 0.25 ;
      LAYER M2 ;
      RECT 408.74 0.0 408.88 0.25 ;
      LAYER M3 ;
      RECT 408.74 0.0 408.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[58]
  PIN DA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 33.55 0.0 33.69 0.25 ;
      LAYER M2 ;
      RECT 33.55 0.0 33.69 0.25 ;
      LAYER M1 ;
      RECT 33.55 0.0 33.69 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[5]
  PIN QA[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 409.525 0.0 409.665 0.25 ;
      LAYER M2 ;
      RECT 409.525 0.0 409.665 0.25 ;
      LAYER M3 ;
      RECT 409.525 0.0 409.665 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[58]
  PIN QA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 32.765 0.0 32.905 0.25 ;
      LAYER M2 ;
      RECT 32.765 0.0 32.905 0.25 ;
      LAYER M1 ;
      RECT 32.765 0.0 32.905 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[5]
  PIN TDA[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 409.905 0.0 410.045 0.25 ;
      LAYER M2 ;
      RECT 409.905 0.0 410.045 0.25 ;
      LAYER M3 ;
      RECT 409.905 0.0 410.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[58]
  PIN TDA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 32.385 0.0 32.525 0.25 ;
      LAYER M2 ;
      RECT 32.385 0.0 32.525 0.25 ;
      LAYER M1 ;
      RECT 32.385 0.0 32.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[5]
  PIN TDB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 410.47 0.0 410.61 0.25 ;
      LAYER M2 ;
      RECT 410.47 0.0 410.61 0.25 ;
      LAYER M3 ;
      RECT 410.47 0.0 410.61 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[59]
  PIN TDB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 31.82 0.0 31.96 0.25 ;
      LAYER M2 ;
      RECT 31.82 0.0 31.96 0.25 ;
      LAYER M1 ;
      RECT 31.82 0.0 31.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[4]
  PIN QB[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 410.855 0.0 410.995 0.25 ;
      LAYER M2 ;
      RECT 410.855 0.0 410.995 0.25 ;
      LAYER M3 ;
      RECT 410.855 0.0 410.995 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[59]
  PIN QB[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 31.435 0.0 31.575 0.25 ;
      LAYER M2 ;
      RECT 31.435 0.0 31.575 0.25 ;
      LAYER M1 ;
      RECT 31.435 0.0 31.575 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[4]
  PIN DB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 411.63 0.0 411.77 0.25 ;
      LAYER M2 ;
      RECT 411.63 0.0 411.77 0.25 ;
      LAYER M3 ;
      RECT 411.63 0.0 411.77 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[59]
  PIN DB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 30.66 0.0 30.8 0.25 ;
      LAYER M2 ;
      RECT 30.66 0.0 30.8 0.25 ;
      LAYER M1 ;
      RECT 30.66 0.0 30.8 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[4]
  PIN DA[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 414.94 0.0 415.08 0.25 ;
      LAYER M2 ;
      RECT 414.94 0.0 415.08 0.25 ;
      LAYER M3 ;
      RECT 414.94 0.0 415.08 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[59]
  PIN DA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 27.35 0.0 27.49 0.25 ;
      LAYER M2 ;
      RECT 27.35 0.0 27.49 0.25 ;
      LAYER M1 ;
      RECT 27.35 0.0 27.49 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[4]
  PIN QA[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 415.725 0.0 415.865 0.25 ;
      LAYER M2 ;
      RECT 415.725 0.0 415.865 0.25 ;
      LAYER M3 ;
      RECT 415.725 0.0 415.865 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[59]
  PIN QA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 26.565 0.0 26.705 0.25 ;
      LAYER M2 ;
      RECT 26.565 0.0 26.705 0.25 ;
      LAYER M1 ;
      RECT 26.565 0.0 26.705 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[4]
  PIN TDA[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 416.105 0.0 416.245 0.25 ;
      LAYER M2 ;
      RECT 416.105 0.0 416.245 0.25 ;
      LAYER M3 ;
      RECT 416.105 0.0 416.245 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[59]
  PIN TDA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 26.185 0.0 26.325 0.25 ;
      LAYER M2 ;
      RECT 26.185 0.0 26.325 0.25 ;
      LAYER M1 ;
      RECT 26.185 0.0 26.325 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[4]
  PIN TDB[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 416.67 0.0 416.81 0.25 ;
      LAYER M2 ;
      RECT 416.67 0.0 416.81 0.25 ;
      LAYER M3 ;
      RECT 416.67 0.0 416.81 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[60]
  PIN TDB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.62 0.0 25.76 0.25 ;
      LAYER M2 ;
      RECT 25.62 0.0 25.76 0.25 ;
      LAYER M1 ;
      RECT 25.62 0.0 25.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[3]
  PIN QB[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 417.055 0.0 417.195 0.25 ;
      LAYER M2 ;
      RECT 417.055 0.0 417.195 0.25 ;
      LAYER M3 ;
      RECT 417.055 0.0 417.195 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[60]
  PIN QB[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.235 0.0 25.375 0.25 ;
      LAYER M2 ;
      RECT 25.235 0.0 25.375 0.25 ;
      LAYER M1 ;
      RECT 25.235 0.0 25.375 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[3]
  PIN DB[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 417.83 0.0 417.97 0.25 ;
      LAYER M2 ;
      RECT 417.83 0.0 417.97 0.25 ;
      LAYER M3 ;
      RECT 417.83 0.0 417.97 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[60]
  PIN DB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 24.46 0.0 24.6 0.25 ;
      LAYER M2 ;
      RECT 24.46 0.0 24.6 0.25 ;
      LAYER M1 ;
      RECT 24.46 0.0 24.6 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[3]
  PIN DA[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 421.14 0.0 421.28 0.25 ;
      LAYER M2 ;
      RECT 421.14 0.0 421.28 0.25 ;
      LAYER M3 ;
      RECT 421.14 0.0 421.28 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[60]
  PIN DA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 21.15 0.0 21.29 0.25 ;
      LAYER M2 ;
      RECT 21.15 0.0 21.29 0.25 ;
      LAYER M1 ;
      RECT 21.15 0.0 21.29 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[3]
  PIN QA[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 421.925 0.0 422.065 0.25 ;
      LAYER M2 ;
      RECT 421.925 0.0 422.065 0.25 ;
      LAYER M3 ;
      RECT 421.925 0.0 422.065 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[60]
  PIN QA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 20.365 0.0 20.505 0.25 ;
      LAYER M2 ;
      RECT 20.365 0.0 20.505 0.25 ;
      LAYER M1 ;
      RECT 20.365 0.0 20.505 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[3]
  PIN TDA[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 422.305 0.0 422.445 0.25 ;
      LAYER M2 ;
      RECT 422.305 0.0 422.445 0.25 ;
      LAYER M3 ;
      RECT 422.305 0.0 422.445 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[60]
  PIN TDA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.985 0.0 20.125 0.25 ;
      LAYER M2 ;
      RECT 19.985 0.0 20.125 0.25 ;
      LAYER M1 ;
      RECT 19.985 0.0 20.125 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[3]
  PIN TDB[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 422.87 0.0 423.01 0.25 ;
      LAYER M2 ;
      RECT 422.87 0.0 423.01 0.25 ;
      LAYER M3 ;
      RECT 422.87 0.0 423.01 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[61]
  PIN TDB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.42 0.0 19.56 0.25 ;
      LAYER M2 ;
      RECT 19.42 0.0 19.56 0.25 ;
      LAYER M1 ;
      RECT 19.42 0.0 19.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[2]
  PIN QB[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 423.255 0.0 423.395 0.25 ;
      LAYER M2 ;
      RECT 423.255 0.0 423.395 0.25 ;
      LAYER M3 ;
      RECT 423.255 0.0 423.395 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[61]
  PIN QB[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.035 0.0 19.175 0.25 ;
      LAYER M2 ;
      RECT 19.035 0.0 19.175 0.25 ;
      LAYER M1 ;
      RECT 19.035 0.0 19.175 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[2]
  PIN DB[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 424.03 0.0 424.17 0.25 ;
      LAYER M2 ;
      RECT 424.03 0.0 424.17 0.25 ;
      LAYER M3 ;
      RECT 424.03 0.0 424.17 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[61]
  PIN DB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 18.26 0.0 18.4 0.25 ;
      LAYER M2 ;
      RECT 18.26 0.0 18.4 0.25 ;
      LAYER M1 ;
      RECT 18.26 0.0 18.4 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[2]
  PIN DA[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 427.34 0.0 427.48 0.25 ;
      LAYER M2 ;
      RECT 427.34 0.0 427.48 0.25 ;
      LAYER M3 ;
      RECT 427.34 0.0 427.48 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[61]
  PIN DA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.95 0.0 15.09 0.25 ;
      LAYER M2 ;
      RECT 14.95 0.0 15.09 0.25 ;
      LAYER M1 ;
      RECT 14.95 0.0 15.09 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[2]
  PIN QA[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 428.125 0.0 428.265 0.25 ;
      LAYER M2 ;
      RECT 428.125 0.0 428.265 0.25 ;
      LAYER M3 ;
      RECT 428.125 0.0 428.265 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[61]
  PIN QA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 14.165 0.0 14.305 0.25 ;
      LAYER M2 ;
      RECT 14.165 0.0 14.305 0.25 ;
      LAYER M1 ;
      RECT 14.165 0.0 14.305 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[2]
  PIN TDA[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 428.505 0.0 428.645 0.25 ;
      LAYER M2 ;
      RECT 428.505 0.0 428.645 0.25 ;
      LAYER M3 ;
      RECT 428.505 0.0 428.645 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[61]
  PIN TDA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.785 0.0 13.925 0.25 ;
      LAYER M2 ;
      RECT 13.785 0.0 13.925 0.25 ;
      LAYER M1 ;
      RECT 13.785 0.0 13.925 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[2]
  PIN TDB[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 429.07 0.0 429.21 0.25 ;
      LAYER M2 ;
      RECT 429.07 0.0 429.21 0.25 ;
      LAYER M3 ;
      RECT 429.07 0.0 429.21 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[62]
  PIN TDB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 13.22 0.0 13.36 0.25 ;
      LAYER M2 ;
      RECT 13.22 0.0 13.36 0.25 ;
      LAYER M1 ;
      RECT 13.22 0.0 13.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[1]
  PIN QB[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 429.455 0.0 429.595 0.25 ;
      LAYER M2 ;
      RECT 429.455 0.0 429.595 0.25 ;
      LAYER M3 ;
      RECT 429.455 0.0 429.595 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[62]
  PIN QB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.835 0.0 12.975 0.25 ;
      LAYER M2 ;
      RECT 12.835 0.0 12.975 0.25 ;
      LAYER M1 ;
      RECT 12.835 0.0 12.975 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[1]
  PIN DB[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 430.23 0.0 430.37 0.25 ;
      LAYER M2 ;
      RECT 430.23 0.0 430.37 0.25 ;
      LAYER M3 ;
      RECT 430.23 0.0 430.37 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[62]
  PIN DB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.06 0.0 12.2 0.25 ;
      LAYER M2 ;
      RECT 12.06 0.0 12.2 0.25 ;
      LAYER M1 ;
      RECT 12.06 0.0 12.2 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[1]
  PIN DA[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 433.54 0.0 433.68 0.25 ;
      LAYER M2 ;
      RECT 433.54 0.0 433.68 0.25 ;
      LAYER M3 ;
      RECT 433.54 0.0 433.68 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[62]
  PIN DA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.75 0.0 8.89 0.25 ;
      LAYER M2 ;
      RECT 8.75 0.0 8.89 0.25 ;
      LAYER M1 ;
      RECT 8.75 0.0 8.89 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[1]
  PIN QA[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 434.325 0.0 434.465 0.25 ;
      LAYER M2 ;
      RECT 434.325 0.0 434.465 0.25 ;
      LAYER M3 ;
      RECT 434.325 0.0 434.465 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[62]
  PIN QA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.965 0.0 8.105 0.25 ;
      LAYER M2 ;
      RECT 7.965 0.0 8.105 0.25 ;
      LAYER M1 ;
      RECT 7.965 0.0 8.105 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[1]
  PIN TDA[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 434.705 0.0 434.845 0.25 ;
      LAYER M2 ;
      RECT 434.705 0.0 434.845 0.25 ;
      LAYER M3 ;
      RECT 434.705 0.0 434.845 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[62]
  PIN TDA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.585 0.0 7.725 0.25 ;
      LAYER M2 ;
      RECT 7.585 0.0 7.725 0.25 ;
      LAYER M1 ;
      RECT 7.585 0.0 7.725 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[1]
  PIN TDB[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 435.27 0.0 435.41 0.25 ;
      LAYER M2 ;
      RECT 435.27 0.0 435.41 0.25 ;
      LAYER M3 ;
      RECT 435.27 0.0 435.41 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[63]
  PIN TDB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.02 0.0 7.16 0.25 ;
      LAYER M2 ;
      RECT 7.02 0.0 7.16 0.25 ;
      LAYER M1 ;
      RECT 7.02 0.0 7.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDB[0]
  PIN QB[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 435.655 0.0 435.795 0.25 ;
      LAYER M2 ;
      RECT 435.655 0.0 435.795 0.25 ;
      LAYER M3 ;
      RECT 435.655 0.0 435.795 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[63]
  PIN QB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.635 0.0 6.775 0.25 ;
      LAYER M2 ;
      RECT 6.635 0.0 6.775 0.25 ;
      LAYER M1 ;
      RECT 6.635 0.0 6.775 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QB[0]
  PIN DB[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 436.43 0.0 436.57 0.25 ;
      LAYER M2 ;
      RECT 436.43 0.0 436.57 0.25 ;
      LAYER M3 ;
      RECT 436.43 0.0 436.57 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[63]
  PIN DB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.86 0.0 6.0 0.25 ;
      LAYER M2 ;
      RECT 5.86 0.0 6.0 0.25 ;
      LAYER M1 ;
      RECT 5.86 0.0 6.0 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[0]
  PIN DA[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 439.74 0.0 439.88 0.25 ;
      LAYER M2 ;
      RECT 439.74 0.0 439.88 0.25 ;
      LAYER M3 ;
      RECT 439.74 0.0 439.88 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[63]
  PIN DA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.55 0.0 2.69 0.25 ;
      LAYER M2 ;
      RECT 2.55 0.0 2.69 0.25 ;
      LAYER M1 ;
      RECT 2.55 0.0 2.69 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DA[0]
  PIN QA[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 440.525 0.0 440.665 0.25 ;
      LAYER M2 ;
      RECT 440.525 0.0 440.665 0.25 ;
      LAYER M3 ;
      RECT 440.525 0.0 440.665 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[63]
  PIN QA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.765 0.0 1.905 0.25 ;
      LAYER M2 ;
      RECT 1.765 0.0 1.905 0.25 ;
      LAYER M1 ;
      RECT 1.765 0.0 1.905 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[0]
  PIN TDA[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 440.905 0.0 441.045 0.25 ;
      LAYER M2 ;
      RECT 440.905 0.0 441.045 0.25 ;
      LAYER M3 ;
      RECT 440.905 0.0 441.045 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[63]
  PIN TDA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.385 0.0 1.525 0.25 ;
      LAYER M2 ;
      RECT 1.385 0.0 1.525 0.25 ;
      LAYER M1 ;
      RECT 1.385 0.0 1.525 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END TDA[0]
  PIN SIA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 441.31 0.0 441.45 0.25 ;
      LAYER M2 ;
      RECT 441.31 0.0 441.45 0.25 ;
      LAYER M3 ;
      RECT 441.31 0.0 441.45 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END SIA[1]
  PIN SIA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.98 0.0 1.12 0.25 ;
      LAYER M2 ;
      RECT 0.98 0.0 1.12 0.25 ;
      LAYER M1 ;
      RECT 0.98 0.0 1.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END SIA[0]
  PIN SIB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 441.87 0.0 442.01 0.25 ;
      LAYER M2 ;
      RECT 441.87 0.0 442.01 0.25 ;
      LAYER M3 ;
      RECT 441.87 0.0 442.01 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END SIB[1]
  PIN SIB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.42 0.0 0.56 0.25 ;
      LAYER M2 ;
      RECT 0.42 0.0 0.56 0.25 ;
      LAYER M1 ;
      RECT 0.42 0.0 0.56 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END SIB[0]
  PIN VDDCE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.605 0.0 2.815 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 5.705 0.0 5.915 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 8.805 0.0 9.015 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 11.905 0.0 12.115 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 15.005 0.0 15.215 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 18.105 0.0 18.315 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 21.205 0.0 21.415 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 24.305 0.0 24.515 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 27.405 0.0 27.615 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 30.505 0.0 30.715 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 33.605 0.0 33.815 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 36.705 0.0 36.915 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 39.805 0.0 40.015 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 42.905 0.0 43.115 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 46.005 0.0 46.215 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 49.105 0.0 49.315 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 52.205 0.0 52.415 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.305 0.0 55.515 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 58.405 0.0 58.615 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 61.505 0.0 61.715 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.605 0.0 64.815 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 67.705 0.0 67.915 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 70.805 0.0 71.015 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 73.905 0.0 74.115 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 77.005 0.0 77.215 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 80.105 0.0 80.315 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 83.205 0.0 83.415 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 86.305 0.0 86.515 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 89.405 0.0 89.615 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 92.505 0.0 92.715 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 95.605 0.0 95.815 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.705 0.0 98.915 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 101.805 0.0 102.015 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 104.905 0.0 105.115 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 108.005 0.0 108.215 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 111.105 0.0 111.315 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 114.205 0.0 114.415 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 117.305 0.0 117.515 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 120.405 0.0 120.615 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 123.505 0.0 123.715 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 126.605 0.0 126.815 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 129.705 0.0 129.915 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 132.805 0.0 133.015 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 135.905 0.0 136.115 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 139.005 0.0 139.215 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 142.105 0.0 142.315 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 145.205 0.0 145.415 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 148.305 0.0 148.515 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 151.405 0.0 151.615 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 154.505 0.0 154.715 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 157.605 0.0 157.815 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 160.705 0.0 160.915 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 163.805 0.0 164.015 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 166.905 0.0 167.115 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 170.005 0.0 170.215 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 173.105 0.0 173.315 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 176.205 0.0 176.415 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 179.305 0.0 179.515 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 182.405 0.0 182.615 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 185.505 0.0 185.715 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 188.605 0.0 188.815 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 191.705 0.0 191.915 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 194.805 0.0 195.015 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 197.905 0.0 198.115 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 204.55 0.0 204.76 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 207.1 0.0 207.31 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 212.215 0.0 212.425 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 212.995 0.0 213.205 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.765 0.0 213.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 214.935 0.0 215.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 216.36 0.0 216.57 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 217.98 0.0 218.19 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 220.21 0.0 220.42 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 222.01 0.0 222.22 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 224.24 0.0 224.45 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 225.86 0.0 226.07 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 227.285 0.0 227.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 228.455 0.0 228.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 229.225 0.0 229.435 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 230.005 0.0 230.215 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 235.12 0.0 235.33 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 237.67 0.0 237.88 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 244.315 0.0 244.525 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 247.415 0.0 247.625 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 250.515 0.0 250.725 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 253.615 0.0 253.825 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 256.715 0.0 256.925 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 259.815 0.0 260.025 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 262.915 0.0 263.125 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 266.015 0.0 266.225 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 269.115 0.0 269.325 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 272.215 0.0 272.425 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 275.315 0.0 275.525 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 278.415 0.0 278.625 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 281.515 0.0 281.725 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 284.615 0.0 284.825 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 287.715 0.0 287.925 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 290.815 0.0 291.025 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 293.915 0.0 294.125 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 297.015 0.0 297.225 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 300.115 0.0 300.325 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 303.215 0.0 303.425 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 306.315 0.0 306.525 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 309.415 0.0 309.625 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 312.515 0.0 312.725 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 315.615 0.0 315.825 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 318.715 0.0 318.925 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 321.815 0.0 322.025 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 324.915 0.0 325.125 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 328.015 0.0 328.225 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 331.115 0.0 331.325 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 334.215 0.0 334.425 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 337.315 0.0 337.525 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 340.415 0.0 340.625 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 343.515 0.0 343.725 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 346.615 0.0 346.825 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 349.715 0.0 349.925 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 352.815 0.0 353.025 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 355.915 0.0 356.125 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 359.015 0.0 359.225 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 362.115 0.0 362.325 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 365.215 0.0 365.425 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 368.315 0.0 368.525 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 371.415 0.0 371.625 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 374.515 0.0 374.725 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 377.615 0.0 377.825 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 380.715 0.0 380.925 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 383.815 0.0 384.025 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 386.915 0.0 387.125 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 390.015 0.0 390.225 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 393.115 0.0 393.325 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 396.215 0.0 396.425 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 399.315 0.0 399.525 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 402.415 0.0 402.625 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 405.515 0.0 405.725 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 408.615 0.0 408.825 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 411.715 0.0 411.925 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 414.815 0.0 415.025 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 417.915 0.0 418.125 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 421.015 0.0 421.225 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 424.115 0.0 424.325 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 427.215 0.0 427.425 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 430.315 0.0 430.525 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 433.415 0.0 433.625 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 436.515 0.0 436.725 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 439.615 0.0 439.825 69.945 ;
      END
    END VDDCE
  PIN VDDPE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 1.055 0.0 1.265 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 4.155 0.0 4.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.255 0.0 7.465 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 10.355 0.0 10.565 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 13.455 0.0 13.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 16.555 0.0 16.765 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 19.655 0.0 19.865 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 22.755 0.0 22.965 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.855 0.0 26.065 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.955 0.0 29.165 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 32.055 0.0 32.265 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.155 0.0 35.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.255 0.0 38.465 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 41.355 0.0 41.565 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.455 0.0 44.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 47.555 0.0 47.765 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 50.655 0.0 50.865 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 53.755 0.0 53.965 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 56.855 0.0 57.065 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 59.955 0.0 60.165 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 63.055 0.0 63.265 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 66.155 0.0 66.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 69.255 0.0 69.465 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.355 0.0 72.565 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 75.455 0.0 75.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 78.555 0.0 78.765 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.655 0.0 81.865 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 84.755 0.0 84.965 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 87.855 0.0 88.065 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 90.955 0.0 91.165 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 94.055 0.0 94.265 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 97.155 0.0 97.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.255 0.0 100.465 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.355 0.0 103.565 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 106.455 0.0 106.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 109.555 0.0 109.765 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 112.655 0.0 112.865 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 115.755 0.0 115.965 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.855 0.0 119.065 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 121.955 0.0 122.165 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 125.055 0.0 125.265 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.155 0.0 128.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 131.255 0.0 131.465 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 134.355 0.0 134.565 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 137.455 0.0 137.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 140.555 0.0 140.765 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 143.655 0.0 143.865 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 146.755 0.0 146.965 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 149.855 0.0 150.065 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 152.955 0.0 153.165 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 156.055 0.0 156.265 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 159.155 0.0 159.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 162.255 0.0 162.465 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 165.355 0.0 165.565 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 168.455 0.0 168.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 171.555 0.0 171.765 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 174.655 0.0 174.865 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 177.755 0.0 177.965 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 180.855 0.0 181.065 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 183.955 0.0 184.165 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 187.055 0.0 187.265 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 190.155 0.0 190.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 193.255 0.0 193.465 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 196.355 0.0 196.565 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 199.455 0.0 199.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 201.985 0.0 202.195 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 202.985 0.0 203.195 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 203.765 0.0 203.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 204.94 0.0 205.15 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 207.88 0.0 208.09 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 211.09 0.0 211.35 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 214.155 0.0 214.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 215.97 0.0 216.18 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 217.18 0.0 217.39 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 218.58 0.0 218.84 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 223.59 0.0 223.85 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 225.04 0.0 225.25 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 226.25 0.0 226.46 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 228.065 0.0 228.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 231.08 0.0 231.34 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 234.34 0.0 234.55 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 237.28 0.0 237.49 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 238.455 0.0 238.665 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 239.235 0.0 239.445 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 240.235 0.0 240.445 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 242.765 0.0 242.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 245.865 0.0 246.075 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 248.965 0.0 249.175 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 252.065 0.0 252.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 255.165 0.0 255.375 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 258.265 0.0 258.475 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 261.365 0.0 261.575 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 264.465 0.0 264.675 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 267.565 0.0 267.775 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 270.665 0.0 270.875 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 273.765 0.0 273.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 276.865 0.0 277.075 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 279.965 0.0 280.175 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 283.065 0.0 283.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 286.165 0.0 286.375 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 289.265 0.0 289.475 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 292.365 0.0 292.575 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 295.465 0.0 295.675 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 298.565 0.0 298.775 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 301.665 0.0 301.875 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 304.765 0.0 304.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 307.865 0.0 308.075 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 310.965 0.0 311.175 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 314.065 0.0 314.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 317.165 0.0 317.375 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 320.265 0.0 320.475 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 323.365 0.0 323.575 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 326.465 0.0 326.675 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 329.565 0.0 329.775 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 332.665 0.0 332.875 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 335.765 0.0 335.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 338.865 0.0 339.075 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 341.965 0.0 342.175 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 345.065 0.0 345.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 348.165 0.0 348.375 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 351.265 0.0 351.475 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 354.365 0.0 354.575 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 357.465 0.0 357.675 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 360.565 0.0 360.775 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 363.665 0.0 363.875 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 366.765 0.0 366.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 369.865 0.0 370.075 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 372.965 0.0 373.175 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 376.065 0.0 376.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 379.165 0.0 379.375 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 382.265 0.0 382.475 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 385.365 0.0 385.575 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 388.465 0.0 388.675 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 391.565 0.0 391.775 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 394.665 0.0 394.875 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 397.765 0.0 397.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 400.865 0.0 401.075 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 403.965 0.0 404.175 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 407.065 0.0 407.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 410.165 0.0 410.375 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 413.265 0.0 413.475 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 416.365 0.0 416.575 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 419.465 0.0 419.675 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 422.565 0.0 422.775 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 425.665 0.0 425.875 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 428.765 0.0 428.975 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 431.865 0.0 432.075 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 434.965 0.0 435.175 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 438.065 0.0 438.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 441.165 0.0 441.375 69.945 ;
      END
    END VDDPE
  PIN VSSE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.625 0.0 1.835 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 4.735 0.0 4.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 6.685 0.0 6.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.825 0.0 8.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 10.935 0.0 11.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 12.885 0.0 13.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 14.025 0.0 14.235 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 17.135 0.0 17.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 19.085 0.0 19.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 20.225 0.0 20.435 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 23.335 0.0 23.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.285 0.0 25.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 26.425 0.0 26.635 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 29.535 0.0 29.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 31.485 0.0 31.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 32.625 0.0 32.835 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.735 0.0 35.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.685 0.0 37.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.825 0.0 39.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 41.935 0.0 42.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 43.885 0.0 44.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.025 0.0 45.235 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 48.135 0.0 48.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 50.085 0.0 50.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 51.225 0.0 51.435 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 54.335 0.0 54.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 56.285 0.0 56.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 57.425 0.0 57.635 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 60.535 0.0 60.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 62.485 0.0 62.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 63.625 0.0 63.835 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 66.735 0.0 66.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 68.685 0.0 68.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 69.825 0.0 70.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.935 0.0 73.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.885 0.0 75.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 76.025 0.0 76.235 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 79.135 0.0 79.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.085 0.0 81.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 82.225 0.0 82.435 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 85.335 0.0 85.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 87.285 0.0 87.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 88.425 0.0 88.635 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 91.535 0.0 91.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 93.485 0.0 93.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 94.625 0.0 94.835 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 97.735 0.0 97.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 99.685 0.0 99.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.825 0.0 101.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.935 0.0 104.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 105.885 0.0 106.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 107.025 0.0 107.235 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 110.135 0.0 110.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 112.085 0.0 112.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 113.225 0.0 113.435 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 116.335 0.0 116.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 118.285 0.0 118.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 119.425 0.0 119.635 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 122.535 0.0 122.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 124.485 0.0 124.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 125.625 0.0 125.835 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 128.735 0.0 128.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 130.685 0.0 130.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 131.825 0.0 132.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 134.935 0.0 135.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 136.885 0.0 137.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 138.025 0.0 138.235 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 141.135 0.0 141.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 143.085 0.0 143.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 144.225 0.0 144.435 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 147.335 0.0 147.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 149.285 0.0 149.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 150.425 0.0 150.635 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 153.535 0.0 153.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 155.485 0.0 155.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 156.625 0.0 156.835 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 159.735 0.0 159.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 161.685 0.0 161.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 162.825 0.0 163.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 165.935 0.0 166.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 167.885 0.0 168.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 169.025 0.0 169.235 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 172.135 0.0 172.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 174.085 0.0 174.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 175.225 0.0 175.435 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 178.335 0.0 178.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 180.285 0.0 180.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 181.425 0.0 181.635 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 184.535 0.0 184.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 186.485 0.0 186.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 187.625 0.0 187.835 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 190.735 0.0 190.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 192.685 0.0 192.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 193.825 0.0 194.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 196.935 0.0 197.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 198.885 0.0 199.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 201.195 0.0 201.405 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 203.375 0.0 203.585 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 204.155 0.0 204.365 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 205.33 0.0 205.54 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 206.57 0.0 206.85 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 207.49 0.0 207.7 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 208.66 0.0 208.87 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 209.825 0.0 210.105 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 211.825 0.0 212.035 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 213.375 0.0 213.585 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 215.585 0.0 215.795 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 220.72 0.0 220.93 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 221.5 0.0 221.71 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 226.635 0.0 226.845 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 228.845 0.0 229.055 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 230.395 0.0 230.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 232.325 0.0 232.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 233.56 0.0 233.77 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 234.73 0.0 234.94 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 235.58 0.0 235.86 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 236.89 0.0 237.1 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 238.065 0.0 238.275 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 238.845 0.0 239.055 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 241.025 0.0 241.235 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 243.335 0.0 243.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 245.285 0.0 245.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 248.395 0.0 248.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 249.535 0.0 249.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 251.485 0.0 251.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 254.595 0.0 254.805 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 255.735 0.0 255.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 257.685 0.0 257.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 260.795 0.0 261.005 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 261.935 0.0 262.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 263.885 0.0 264.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 266.995 0.0 267.205 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 268.135 0.0 268.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 270.085 0.0 270.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 273.195 0.0 273.405 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 274.335 0.0 274.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 276.285 0.0 276.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 279.395 0.0 279.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 280.535 0.0 280.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 282.485 0.0 282.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 285.595 0.0 285.805 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 286.735 0.0 286.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 288.685 0.0 288.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 291.795 0.0 292.005 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 292.935 0.0 293.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 294.885 0.0 295.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 297.995 0.0 298.205 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 299.135 0.0 299.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 301.085 0.0 301.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 304.195 0.0 304.405 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 305.335 0.0 305.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 307.285 0.0 307.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 310.395 0.0 310.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 311.535 0.0 311.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 313.485 0.0 313.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 316.595 0.0 316.805 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 317.735 0.0 317.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 319.685 0.0 319.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 322.795 0.0 323.005 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 323.935 0.0 324.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 325.885 0.0 326.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 328.995 0.0 329.205 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 330.135 0.0 330.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 332.085 0.0 332.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 335.195 0.0 335.405 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 336.335 0.0 336.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 338.285 0.0 338.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 341.395 0.0 341.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 342.535 0.0 342.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 344.485 0.0 344.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 347.595 0.0 347.805 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 348.735 0.0 348.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 350.685 0.0 350.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 353.795 0.0 354.005 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 354.935 0.0 355.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 356.885 0.0 357.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 359.995 0.0 360.205 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 361.135 0.0 361.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 363.085 0.0 363.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 366.195 0.0 366.405 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 367.335 0.0 367.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 369.285 0.0 369.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 372.395 0.0 372.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 373.535 0.0 373.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 375.485 0.0 375.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 378.595 0.0 378.805 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 379.735 0.0 379.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 381.685 0.0 381.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 384.795 0.0 385.005 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 385.935 0.0 386.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 387.885 0.0 388.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 390.995 0.0 391.205 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 392.135 0.0 392.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 394.085 0.0 394.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 397.195 0.0 397.405 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 398.335 0.0 398.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 400.285 0.0 400.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 403.395 0.0 403.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 404.535 0.0 404.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 406.485 0.0 406.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 409.595 0.0 409.805 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 410.735 0.0 410.945 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 412.685 0.0 412.895 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 415.795 0.0 416.005 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 416.935 0.0 417.145 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 418.885 0.0 419.095 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 421.995 0.0 422.205 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 423.135 0.0 423.345 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 425.085 0.0 425.295 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 428.195 0.0 428.405 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 429.335 0.0 429.545 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 431.285 0.0 431.495 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 434.395 0.0 434.605 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 435.535 0.0 435.745 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 437.485 0.0 437.695 69.945 ;
      END
    PORT
      LAYER M4 ;
      RECT 440.595 0.0 440.805 69.945 ;
      END
    END VSSE
  OBS
    #otc obstructions
    LAYER M1 DESIGNRULEWIDTH 0.07 ;
    RECT 442.15 0.0 442.43 0.32 ;
    RECT 441.59 0.0 441.73 0.32 ;
    RECT 440.02 0.0 440.385 0.32 ;
    RECT 436.71 0.0 439.6 0.32 ;
    RECT 435.935 0.0 436.29 0.32 ;
    RECT 434.985 0.0 435.13 0.32 ;
    RECT 433.82 0.0 434.185 0.32 ;
    RECT 430.51 0.0 433.4 0.32 ;
    RECT 429.735 0.0 430.09 0.32 ;
    RECT 428.785 0.0 428.93 0.32 ;
    RECT 427.62 0.0 427.985 0.32 ;
    RECT 424.31 0.0 427.2 0.32 ;
    RECT 423.535 0.0 423.89 0.32 ;
    RECT 422.585 0.0 422.73 0.32 ;
    RECT 421.42 0.0 421.785 0.32 ;
    RECT 418.11 0.0 421.0 0.32 ;
    RECT 417.335 0.0 417.69 0.32 ;
    RECT 416.385 0.0 416.53 0.32 ;
    RECT 415.22 0.0 415.585 0.32 ;
    RECT 411.91 0.0 414.8 0.32 ;
    RECT 411.135 0.0 411.49 0.32 ;
    RECT 410.185 0.0 410.33 0.32 ;
    RECT 409.02 0.0 409.385 0.32 ;
    RECT 405.71 0.0 408.6 0.32 ;
    RECT 404.935 0.0 405.29 0.32 ;
    RECT 403.985 0.0 404.13 0.32 ;
    RECT 402.82 0.0 403.185 0.32 ;
    RECT 399.51 0.0 402.4 0.32 ;
    RECT 398.735 0.0 399.09 0.32 ;
    RECT 397.785 0.0 397.93 0.32 ;
    RECT 396.62 0.0 396.985 0.32 ;
    RECT 393.31 0.0 396.2 0.32 ;
    RECT 392.535 0.0 392.89 0.32 ;
    RECT 391.585 0.0 391.73 0.32 ;
    RECT 390.42 0.0 390.785 0.32 ;
    RECT 387.11 0.0 390.0 0.32 ;
    RECT 386.335 0.0 386.69 0.32 ;
    RECT 385.385 0.0 385.53 0.32 ;
    RECT 384.22 0.0 384.585 0.32 ;
    RECT 380.91 0.0 383.8 0.32 ;
    RECT 380.135 0.0 380.49 0.32 ;
    RECT 379.185 0.0 379.33 0.32 ;
    RECT 378.02 0.0 378.385 0.32 ;
    RECT 374.71 0.0 377.6 0.32 ;
    RECT 373.935 0.0 374.29 0.32 ;
    RECT 372.985 0.0 373.13 0.32 ;
    RECT 371.82 0.0 372.185 0.32 ;
    RECT 368.51 0.0 371.4 0.32 ;
    RECT 367.735 0.0 368.09 0.32 ;
    RECT 366.785 0.0 366.93 0.32 ;
    RECT 365.62 0.0 365.985 0.32 ;
    RECT 362.31 0.0 365.2 0.32 ;
    RECT 361.535 0.0 361.89 0.32 ;
    RECT 360.585 0.0 360.73 0.32 ;
    RECT 359.42 0.0 359.785 0.32 ;
    RECT 356.11 0.0 359.0 0.32 ;
    RECT 355.335 0.0 355.69 0.32 ;
    RECT 354.385 0.0 354.53 0.32 ;
    RECT 353.22 0.0 353.585 0.32 ;
    RECT 349.91 0.0 352.8 0.32 ;
    RECT 349.135 0.0 349.49 0.32 ;
    RECT 348.185 0.0 348.33 0.32 ;
    RECT 347.02 0.0 347.385 0.32 ;
    RECT 343.71 0.0 346.6 0.32 ;
    RECT 342.935 0.0 343.29 0.32 ;
    RECT 341.985 0.0 342.13 0.32 ;
    RECT 340.82 0.0 341.185 0.32 ;
    RECT 337.51 0.0 340.4 0.32 ;
    RECT 336.735 0.0 337.09 0.32 ;
    RECT 335.785 0.0 335.93 0.32 ;
    RECT 334.62 0.0 334.985 0.32 ;
    RECT 331.31 0.0 334.2 0.32 ;
    RECT 330.535 0.0 330.89 0.32 ;
    RECT 329.585 0.0 329.73 0.32 ;
    RECT 328.42 0.0 328.785 0.32 ;
    RECT 325.11 0.0 328.0 0.32 ;
    RECT 324.335 0.0 324.69 0.32 ;
    RECT 323.385 0.0 323.53 0.32 ;
    RECT 322.22 0.0 322.585 0.32 ;
    RECT 318.91 0.0 321.8 0.32 ;
    RECT 318.135 0.0 318.49 0.32 ;
    RECT 317.185 0.0 317.33 0.32 ;
    RECT 316.02 0.0 316.385 0.32 ;
    RECT 312.71 0.0 315.6 0.32 ;
    RECT 311.935 0.0 312.29 0.32 ;
    RECT 310.985 0.0 311.13 0.32 ;
    RECT 309.82 0.0 310.185 0.32 ;
    RECT 306.51 0.0 309.4 0.32 ;
    RECT 305.735 0.0 306.09 0.32 ;
    RECT 304.785 0.0 304.93 0.32 ;
    RECT 303.62 0.0 303.985 0.32 ;
    RECT 300.31 0.0 303.2 0.32 ;
    RECT 299.535 0.0 299.89 0.32 ;
    RECT 298.585 0.0 298.73 0.32 ;
    RECT 297.42 0.0 297.785 0.32 ;
    RECT 294.11 0.0 297.0 0.32 ;
    RECT 293.335 0.0 293.69 0.32 ;
    RECT 291.53 0.0 291.795 0.32 ;
    RECT 290.27 0.0 290.765 0.32 ;
    RECT 289.485 0.0 289.85 0.32 ;
    RECT 287.905 0.0 288.435 0.32 ;
    RECT 286.775 0.0 287.485 0.32 ;
    RECT 286.215 0.0 286.355 0.32 ;
    RECT 285.225 0.0 285.795 0.32 ;
    RECT 281.535 0.0 284.805 0.32 ;
    RECT 280.69 0.0 281.115 0.32 ;
    RECT 280.125 0.0 280.27 0.32 ;
    RECT 279.065 0.0 279.705 0.32 ;
    RECT 276.665 0.0 278.645 0.32 ;
    RECT 275.595 0.0 276.245 0.32 ;
    RECT 274.65 0.0 274.895 0.32 ;
    RECT 273.8 0.0 273.95 0.32 ;
    RECT 272.825 0.0 273.38 0.32 ;
    RECT 271.605 0.0 272.405 0.32 ;
    RECT 270.635 0.0 270.905 0.32 ;
    RECT 269.135 0.0 270.215 0.32 ;
    RECT 268.355 0.0 268.715 0.32 ;
    RECT 266.625 0.0 266.81 0.32 ;
    RECT 263.105 0.0 266.205 0.32 ;
    RECT 262.015 0.0 262.405 0.32 ;
    RECT 260.425 0.0 260.7 0.32 ;
    RECT 257.875 0.0 259.705 0.32 ;
    RECT 257.025 0.0 257.455 0.32 ;
    RECT 256.065 0.0 256.315 0.32 ;
    RECT 255.215 0.0 255.365 0.32 ;
    RECT 254.225 0.0 254.795 0.32 ;
    RECT 253.16 0.0 253.805 0.32 ;
    RECT 252.1 0.0 252.445 0.32 ;
    RECT 250.575 0.0 251.38 0.32 ;
    RECT 249.66 0.0 250.155 0.32 ;
    RECT 249.095 0.0 249.24 0.32 ;
    RECT 248.025 0.0 248.675 0.32 ;
    RECT 244.315 0.0 247.605 0.32 ;
    RECT 243.665 0.0 243.895 0.32 ;
    RECT 241.54 0.0 242.565 0.32 ;
    RECT 240.985 0.0 241.12 0.32 ;
    RECT 239.93 0.0 240.13 0.32 ;
    RECT 238.05 0.0 239.13 0.32 ;
    RECT 235.96 0.0 237.22 0.32 ;
    RECT 231.965 0.0 235.095 0.32 ;
    RECT 231.3 0.0 231.545 0.32 ;
    RECT 230.135 0.0 230.46 0.32 ;
    RECT 222.235 0.0 229.715 0.32 ;
    RECT 211.79 0.0 221.815 0.32 ;
    RECT 210.885 0.0 211.07 0.32 ;
    RECT 207.31 0.0 210.465 0.32 ;
    RECT 206.57 0.0 206.89 0.32 ;
    RECT 205.845 0.0 206.15 0.32 ;
    RECT 203.3 0.0 205.12 0.32 ;
    RECT 202.105 0.0 202.5 0.32 ;
    RECT 201.505 0.0 201.685 0.32 ;
    RECT 200.08 0.0 200.635 0.32 ;
    RECT 199.465 0.0 199.66 0.32 ;
    RECT 198.555 0.0 198.765 0.32 ;
    RECT 194.825 0.0 198.135 0.32 ;
    RECT 193.965 0.0 194.405 0.32 ;
    RECT 193.405 0.0 193.545 0.32 ;
    RECT 192.315 0.0 192.985 0.32 ;
    RECT 190.785 0.0 191.895 0.32 ;
    RECT 188.625 0.0 189.39 0.32 ;
    RECT 187.62 0.0 188.205 0.32 ;
    RECT 186.2 0.0 186.445 0.32 ;
    RECT 184.91 0.0 185.5 0.32 ;
    RECT 182.66 0.0 184.49 0.32 ;
    RECT 181.715 0.0 181.96 0.32 ;
    RECT 179.865 0.0 180.12 0.32 ;
    RECT 176.225 0.0 179.135 0.32 ;
    RECT 175.645 0.0 175.805 0.32 ;
    RECT 173.715 0.0 174.035 0.32 ;
    RECT 171.99 0.0 173.295 0.32 ;
    RECT 171.445 0.0 171.57 0.32 ;
    RECT 170.025 0.0 170.725 0.32 ;
    RECT 169.075 0.0 169.605 0.32 ;
    RECT 168.505 0.0 168.655 0.32 ;
    RECT 167.565 0.0 167.75 0.32 ;
    RECT 166.215 0.0 166.835 0.32 ;
    RECT 163.775 0.0 165.795 0.32 ;
    RECT 162.895 0.0 163.355 0.32 ;
    RECT 162.305 0.0 162.475 0.32 ;
    RECT 161.315 0.0 161.885 0.32 ;
    RECT 157.625 0.0 160.895 0.32 ;
    RECT 156.855 0.0 157.205 0.32 ;
    RECT 156.275 0.0 156.435 0.32 ;
    RECT 155.04 0.0 155.855 0.32 ;
    RECT 154.105 0.0 154.62 0.32 ;
    RECT 152.65 0.0 153.0 0.32 ;
    RECT 151.72 0.0 152.23 0.32 ;
    RECT 150.735 0.0 150.99 0.32 ;
    RECT 149.9 0.0 150.035 0.32 ;
    RECT 148.74 0.0 149.095 0.32 ;
    RECT 145.43 0.0 148.32 0.32 ;
    RECT 144.645 0.0 145.01 0.32 ;
    RECT 143.7 0.0 143.845 0.32 ;
    RECT 142.54 0.0 142.895 0.32 ;
    RECT 139.23 0.0 142.12 0.32 ;
    RECT 138.445 0.0 138.81 0.32 ;
    RECT 137.5 0.0 137.645 0.32 ;
    RECT 136.34 0.0 136.695 0.32 ;
    RECT 133.03 0.0 135.92 0.32 ;
    RECT 132.245 0.0 132.61 0.32 ;
    RECT 131.3 0.0 131.445 0.32 ;
    RECT 130.14 0.0 130.495 0.32 ;
    RECT 126.83 0.0 129.72 0.32 ;
    RECT 126.045 0.0 126.41 0.32 ;
    RECT 125.1 0.0 125.245 0.32 ;
    RECT 123.94 0.0 124.295 0.32 ;
    RECT 120.63 0.0 123.52 0.32 ;
    RECT 119.845 0.0 120.21 0.32 ;
    RECT 118.9 0.0 119.045 0.32 ;
    RECT 117.74 0.0 118.095 0.32 ;
    RECT 114.43 0.0 117.32 0.32 ;
    RECT 113.645 0.0 114.01 0.32 ;
    RECT 112.7 0.0 112.845 0.32 ;
    RECT 111.54 0.0 111.895 0.32 ;
    RECT 108.23 0.0 111.12 0.32 ;
    RECT 107.445 0.0 107.81 0.32 ;
    RECT 106.5 0.0 106.645 0.32 ;
    RECT 105.34 0.0 105.695 0.32 ;
    RECT 102.03 0.0 104.92 0.32 ;
    RECT 101.245 0.0 101.61 0.32 ;
    RECT 100.3 0.0 100.445 0.32 ;
    RECT 99.14 0.0 99.495 0.32 ;
    RECT 95.83 0.0 98.72 0.32 ;
    RECT 95.045 0.0 95.41 0.32 ;
    RECT 94.1 0.0 94.245 0.32 ;
    RECT 92.94 0.0 93.295 0.32 ;
    RECT 89.63 0.0 92.52 0.32 ;
    RECT 88.845 0.0 89.21 0.32 ;
    RECT 87.9 0.0 88.045 0.32 ;
    RECT 86.74 0.0 87.095 0.32 ;
    RECT 83.43 0.0 86.32 0.32 ;
    RECT 82.645 0.0 83.01 0.32 ;
    RECT 81.7 0.0 81.845 0.32 ;
    RECT 80.54 0.0 80.895 0.32 ;
    RECT 77.23 0.0 80.12 0.32 ;
    RECT 76.445 0.0 76.81 0.32 ;
    RECT 75.5 0.0 75.645 0.32 ;
    RECT 74.34 0.0 74.695 0.32 ;
    RECT 71.03 0.0 73.92 0.32 ;
    RECT 70.245 0.0 70.61 0.32 ;
    RECT 69.3 0.0 69.445 0.32 ;
    RECT 68.14 0.0 68.495 0.32 ;
    RECT 64.83 0.0 67.72 0.32 ;
    RECT 64.045 0.0 64.41 0.32 ;
    RECT 63.1 0.0 63.245 0.32 ;
    RECT 61.94 0.0 62.295 0.32 ;
    RECT 58.63 0.0 61.52 0.32 ;
    RECT 57.845 0.0 58.21 0.32 ;
    RECT 56.9 0.0 57.045 0.32 ;
    RECT 55.74 0.0 56.095 0.32 ;
    RECT 52.43 0.0 55.32 0.32 ;
    RECT 51.645 0.0 52.01 0.32 ;
    RECT 50.7 0.0 50.845 0.32 ;
    RECT 49.54 0.0 49.895 0.32 ;
    RECT 46.23 0.0 49.12 0.32 ;
    RECT 45.445 0.0 45.81 0.32 ;
    RECT 44.5 0.0 44.645 0.32 ;
    RECT 43.34 0.0 43.695 0.32 ;
    RECT 40.03 0.0 42.92 0.32 ;
    RECT 39.245 0.0 39.61 0.32 ;
    RECT 38.3 0.0 38.445 0.32 ;
    RECT 37.14 0.0 37.495 0.32 ;
    RECT 33.83 0.0 36.72 0.32 ;
    RECT 33.045 0.0 33.41 0.32 ;
    RECT 32.1 0.0 32.245 0.32 ;
    RECT 30.94 0.0 31.295 0.32 ;
    RECT 27.63 0.0 30.52 0.32 ;
    RECT 26.845 0.0 27.21 0.32 ;
    RECT 25.9 0.0 26.045 0.32 ;
    RECT 24.74 0.0 25.095 0.32 ;
    RECT 21.43 0.0 24.32 0.32 ;
    RECT 20.645 0.0 21.01 0.32 ;
    RECT 19.7 0.0 19.845 0.32 ;
    RECT 18.54 0.0 18.895 0.32 ;
    RECT 15.23 0.0 18.12 0.32 ;
    RECT 14.445 0.0 14.81 0.32 ;
    RECT 13.5 0.0 13.645 0.32 ;
    RECT 12.34 0.0 12.695 0.32 ;
    RECT 9.03 0.0 11.92 0.32 ;
    RECT 8.245 0.0 8.61 0.32 ;
    RECT 7.3 0.0 7.445 0.32 ;
    RECT 6.14 0.0 6.495 0.32 ;
    RECT 2.83 0.0 5.72 0.32 ;
    RECT 2.045 0.0 2.41 0.32 ;
    RECT 0.7 0.0 0.84 0.32 ;
    RECT 0.0 0.0 0.28 0.32 ;
    RECT 0.0 0.32 442.43 69.945 ;
    LAYER V1 ;
    RECT 0.0 0.0 442.43 69.945 ;
    LAYER M2 DESIGNRULEWIDTH 0.07 ;
    RECT 442.15 0.0 442.43 0.32 ;
    RECT 441.59 0.0 441.73 0.32 ;
    RECT 440.02 0.0 440.385 0.32 ;
    RECT 436.71 0.0 439.6 0.32 ;
    RECT 435.935 0.0 436.29 0.32 ;
    RECT 434.985 0.0 435.13 0.32 ;
    RECT 433.82 0.0 434.185 0.32 ;
    RECT 430.51 0.0 433.4 0.32 ;
    RECT 429.735 0.0 430.09 0.32 ;
    RECT 428.785 0.0 428.93 0.32 ;
    RECT 427.62 0.0 427.985 0.32 ;
    RECT 424.31 0.0 427.2 0.32 ;
    RECT 423.535 0.0 423.89 0.32 ;
    RECT 422.585 0.0 422.73 0.32 ;
    RECT 421.42 0.0 421.785 0.32 ;
    RECT 418.11 0.0 421.0 0.32 ;
    RECT 417.335 0.0 417.69 0.32 ;
    RECT 416.385 0.0 416.53 0.32 ;
    RECT 415.22 0.0 415.585 0.32 ;
    RECT 411.91 0.0 414.8 0.32 ;
    RECT 411.135 0.0 411.49 0.32 ;
    RECT 410.185 0.0 410.33 0.32 ;
    RECT 409.02 0.0 409.385 0.32 ;
    RECT 405.71 0.0 408.6 0.32 ;
    RECT 404.935 0.0 405.29 0.32 ;
    RECT 403.985 0.0 404.13 0.32 ;
    RECT 402.82 0.0 403.185 0.32 ;
    RECT 399.51 0.0 402.4 0.32 ;
    RECT 398.735 0.0 399.09 0.32 ;
    RECT 397.785 0.0 397.93 0.32 ;
    RECT 396.62 0.0 396.985 0.32 ;
    RECT 393.31 0.0 396.2 0.32 ;
    RECT 392.535 0.0 392.89 0.32 ;
    RECT 391.585 0.0 391.73 0.32 ;
    RECT 390.42 0.0 390.785 0.32 ;
    RECT 387.11 0.0 390.0 0.32 ;
    RECT 386.335 0.0 386.69 0.32 ;
    RECT 385.385 0.0 385.53 0.32 ;
    RECT 384.22 0.0 384.585 0.32 ;
    RECT 380.91 0.0 383.8 0.32 ;
    RECT 380.135 0.0 380.49 0.32 ;
    RECT 379.185 0.0 379.33 0.32 ;
    RECT 378.02 0.0 378.385 0.32 ;
    RECT 374.71 0.0 377.6 0.32 ;
    RECT 373.935 0.0 374.29 0.32 ;
    RECT 372.985 0.0 373.13 0.32 ;
    RECT 371.82 0.0 372.185 0.32 ;
    RECT 368.51 0.0 371.4 0.32 ;
    RECT 367.735 0.0 368.09 0.32 ;
    RECT 366.785 0.0 366.93 0.32 ;
    RECT 365.62 0.0 365.985 0.32 ;
    RECT 362.31 0.0 365.2 0.32 ;
    RECT 361.535 0.0 361.89 0.32 ;
    RECT 360.585 0.0 360.73 0.32 ;
    RECT 359.42 0.0 359.785 0.32 ;
    RECT 356.11 0.0 359.0 0.32 ;
    RECT 355.335 0.0 355.69 0.32 ;
    RECT 354.385 0.0 354.53 0.32 ;
    RECT 353.22 0.0 353.585 0.32 ;
    RECT 349.91 0.0 352.8 0.32 ;
    RECT 349.135 0.0 349.49 0.32 ;
    RECT 348.185 0.0 348.33 0.32 ;
    RECT 347.02 0.0 347.385 0.32 ;
    RECT 343.71 0.0 346.6 0.32 ;
    RECT 342.935 0.0 343.29 0.32 ;
    RECT 341.985 0.0 342.13 0.32 ;
    RECT 340.82 0.0 341.185 0.32 ;
    RECT 337.51 0.0 340.4 0.32 ;
    RECT 336.735 0.0 337.09 0.32 ;
    RECT 335.785 0.0 335.93 0.32 ;
    RECT 334.62 0.0 334.985 0.32 ;
    RECT 331.31 0.0 334.2 0.32 ;
    RECT 330.535 0.0 330.89 0.32 ;
    RECT 329.585 0.0 329.73 0.32 ;
    RECT 328.42 0.0 328.785 0.32 ;
    RECT 325.11 0.0 328.0 0.32 ;
    RECT 324.335 0.0 324.69 0.32 ;
    RECT 323.385 0.0 323.53 0.32 ;
    RECT 322.22 0.0 322.585 0.32 ;
    RECT 318.91 0.0 321.8 0.32 ;
    RECT 318.135 0.0 318.49 0.32 ;
    RECT 317.185 0.0 317.33 0.32 ;
    RECT 316.02 0.0 316.385 0.32 ;
    RECT 312.71 0.0 315.6 0.32 ;
    RECT 311.935 0.0 312.29 0.32 ;
    RECT 310.985 0.0 311.13 0.32 ;
    RECT 309.82 0.0 310.185 0.32 ;
    RECT 306.51 0.0 309.4 0.32 ;
    RECT 305.735 0.0 306.09 0.32 ;
    RECT 304.785 0.0 304.93 0.32 ;
    RECT 303.62 0.0 303.985 0.32 ;
    RECT 300.31 0.0 303.2 0.32 ;
    RECT 299.535 0.0 299.89 0.32 ;
    RECT 298.585 0.0 298.73 0.32 ;
    RECT 297.42 0.0 297.785 0.32 ;
    RECT 294.11 0.0 297.0 0.32 ;
    RECT 293.335 0.0 293.69 0.32 ;
    RECT 291.53 0.0 291.795 0.32 ;
    RECT 290.27 0.0 290.765 0.32 ;
    RECT 289.485 0.0 289.85 0.32 ;
    RECT 287.905 0.0 288.435 0.32 ;
    RECT 286.775 0.0 287.485 0.32 ;
    RECT 286.215 0.0 286.355 0.32 ;
    RECT 285.225 0.0 285.795 0.32 ;
    RECT 281.535 0.0 284.805 0.32 ;
    RECT 280.69 0.0 281.115 0.32 ;
    RECT 280.125 0.0 280.27 0.32 ;
    RECT 279.065 0.0 279.705 0.32 ;
    RECT 276.665 0.0 278.645 0.32 ;
    RECT 275.595 0.0 276.245 0.32 ;
    RECT 274.65 0.0 274.895 0.32 ;
    RECT 273.8 0.0 273.95 0.32 ;
    RECT 272.825 0.0 273.38 0.32 ;
    RECT 271.605 0.0 272.405 0.32 ;
    RECT 270.635 0.0 270.905 0.32 ;
    RECT 269.135 0.0 270.215 0.32 ;
    RECT 268.355 0.0 268.715 0.32 ;
    RECT 266.625 0.0 266.81 0.32 ;
    RECT 263.105 0.0 266.205 0.32 ;
    RECT 262.015 0.0 262.405 0.32 ;
    RECT 260.425 0.0 260.7 0.32 ;
    RECT 257.875 0.0 259.705 0.32 ;
    RECT 257.025 0.0 257.455 0.32 ;
    RECT 256.065 0.0 256.315 0.32 ;
    RECT 255.215 0.0 255.365 0.32 ;
    RECT 254.225 0.0 254.795 0.32 ;
    RECT 253.16 0.0 253.805 0.32 ;
    RECT 252.1 0.0 252.445 0.32 ;
    RECT 250.575 0.0 251.38 0.32 ;
    RECT 249.66 0.0 250.155 0.32 ;
    RECT 249.095 0.0 249.24 0.32 ;
    RECT 248.025 0.0 248.675 0.32 ;
    RECT 244.315 0.0 247.605 0.32 ;
    RECT 243.665 0.0 243.895 0.32 ;
    RECT 241.54 0.0 242.565 0.32 ;
    RECT 240.985 0.0 241.12 0.32 ;
    RECT 239.93 0.0 240.13 0.32 ;
    RECT 238.05 0.0 239.13 0.32 ;
    RECT 235.96 0.0 237.22 0.32 ;
    RECT 231.965 0.0 235.095 0.32 ;
    RECT 231.3 0.0 231.545 0.32 ;
    RECT 230.135 0.0 230.46 0.32 ;
    RECT 222.235 0.0 229.715 0.32 ;
    RECT 211.79 0.0 221.815 0.32 ;
    RECT 210.885 0.0 211.07 0.32 ;
    RECT 207.31 0.0 210.465 0.32 ;
    RECT 206.57 0.0 206.89 0.32 ;
    RECT 205.845 0.0 206.15 0.32 ;
    RECT 203.3 0.0 205.12 0.32 ;
    RECT 202.105 0.0 202.5 0.32 ;
    RECT 201.505 0.0 201.685 0.32 ;
    RECT 200.08 0.0 200.635 0.32 ;
    RECT 199.465 0.0 199.66 0.32 ;
    RECT 198.555 0.0 198.765 0.32 ;
    RECT 194.825 0.0 198.135 0.32 ;
    RECT 193.965 0.0 194.405 0.32 ;
    RECT 193.405 0.0 193.545 0.32 ;
    RECT 192.315 0.0 192.985 0.32 ;
    RECT 190.785 0.0 191.895 0.32 ;
    RECT 188.625 0.0 189.39 0.32 ;
    RECT 187.62 0.0 188.205 0.32 ;
    RECT 186.2 0.0 186.445 0.32 ;
    RECT 184.91 0.0 185.5 0.32 ;
    RECT 182.66 0.0 184.49 0.32 ;
    RECT 181.715 0.0 181.96 0.32 ;
    RECT 179.865 0.0 180.12 0.32 ;
    RECT 176.225 0.0 179.135 0.32 ;
    RECT 175.645 0.0 175.805 0.32 ;
    RECT 173.715 0.0 174.035 0.32 ;
    RECT 171.99 0.0 173.295 0.32 ;
    RECT 171.445 0.0 171.57 0.32 ;
    RECT 170.025 0.0 170.725 0.32 ;
    RECT 169.075 0.0 169.605 0.32 ;
    RECT 168.505 0.0 168.655 0.32 ;
    RECT 167.565 0.0 167.75 0.32 ;
    RECT 166.215 0.0 166.835 0.32 ;
    RECT 163.775 0.0 165.795 0.32 ;
    RECT 162.895 0.0 163.355 0.32 ;
    RECT 162.305 0.0 162.475 0.32 ;
    RECT 161.315 0.0 161.885 0.32 ;
    RECT 157.625 0.0 160.895 0.32 ;
    RECT 156.855 0.0 157.205 0.32 ;
    RECT 156.275 0.0 156.435 0.32 ;
    RECT 155.04 0.0 155.855 0.32 ;
    RECT 154.105 0.0 154.62 0.32 ;
    RECT 152.65 0.0 153.0 0.32 ;
    RECT 151.72 0.0 152.23 0.32 ;
    RECT 150.735 0.0 150.99 0.32 ;
    RECT 149.9 0.0 150.035 0.32 ;
    RECT 148.74 0.0 149.095 0.32 ;
    RECT 145.43 0.0 148.32 0.32 ;
    RECT 144.645 0.0 145.01 0.32 ;
    RECT 143.7 0.0 143.845 0.32 ;
    RECT 142.54 0.0 142.895 0.32 ;
    RECT 139.23 0.0 142.12 0.32 ;
    RECT 138.445 0.0 138.81 0.32 ;
    RECT 137.5 0.0 137.645 0.32 ;
    RECT 136.34 0.0 136.695 0.32 ;
    RECT 133.03 0.0 135.92 0.32 ;
    RECT 132.245 0.0 132.61 0.32 ;
    RECT 131.3 0.0 131.445 0.32 ;
    RECT 130.14 0.0 130.495 0.32 ;
    RECT 126.83 0.0 129.72 0.32 ;
    RECT 126.045 0.0 126.41 0.32 ;
    RECT 125.1 0.0 125.245 0.32 ;
    RECT 123.94 0.0 124.295 0.32 ;
    RECT 120.63 0.0 123.52 0.32 ;
    RECT 119.845 0.0 120.21 0.32 ;
    RECT 118.9 0.0 119.045 0.32 ;
    RECT 117.74 0.0 118.095 0.32 ;
    RECT 114.43 0.0 117.32 0.32 ;
    RECT 113.645 0.0 114.01 0.32 ;
    RECT 112.7 0.0 112.845 0.32 ;
    RECT 111.54 0.0 111.895 0.32 ;
    RECT 108.23 0.0 111.12 0.32 ;
    RECT 107.445 0.0 107.81 0.32 ;
    RECT 106.5 0.0 106.645 0.32 ;
    RECT 105.34 0.0 105.695 0.32 ;
    RECT 102.03 0.0 104.92 0.32 ;
    RECT 101.245 0.0 101.61 0.32 ;
    RECT 100.3 0.0 100.445 0.32 ;
    RECT 99.14 0.0 99.495 0.32 ;
    RECT 95.83 0.0 98.72 0.32 ;
    RECT 95.045 0.0 95.41 0.32 ;
    RECT 94.1 0.0 94.245 0.32 ;
    RECT 92.94 0.0 93.295 0.32 ;
    RECT 89.63 0.0 92.52 0.32 ;
    RECT 88.845 0.0 89.21 0.32 ;
    RECT 87.9 0.0 88.045 0.32 ;
    RECT 86.74 0.0 87.095 0.32 ;
    RECT 83.43 0.0 86.32 0.32 ;
    RECT 82.645 0.0 83.01 0.32 ;
    RECT 81.7 0.0 81.845 0.32 ;
    RECT 80.54 0.0 80.895 0.32 ;
    RECT 77.23 0.0 80.12 0.32 ;
    RECT 76.445 0.0 76.81 0.32 ;
    RECT 75.5 0.0 75.645 0.32 ;
    RECT 74.34 0.0 74.695 0.32 ;
    RECT 71.03 0.0 73.92 0.32 ;
    RECT 70.245 0.0 70.61 0.32 ;
    RECT 69.3 0.0 69.445 0.32 ;
    RECT 68.14 0.0 68.495 0.32 ;
    RECT 64.83 0.0 67.72 0.32 ;
    RECT 64.045 0.0 64.41 0.32 ;
    RECT 63.1 0.0 63.245 0.32 ;
    RECT 61.94 0.0 62.295 0.32 ;
    RECT 58.63 0.0 61.52 0.32 ;
    RECT 57.845 0.0 58.21 0.32 ;
    RECT 56.9 0.0 57.045 0.32 ;
    RECT 55.74 0.0 56.095 0.32 ;
    RECT 52.43 0.0 55.32 0.32 ;
    RECT 51.645 0.0 52.01 0.32 ;
    RECT 50.7 0.0 50.845 0.32 ;
    RECT 49.54 0.0 49.895 0.32 ;
    RECT 46.23 0.0 49.12 0.32 ;
    RECT 45.445 0.0 45.81 0.32 ;
    RECT 44.5 0.0 44.645 0.32 ;
    RECT 43.34 0.0 43.695 0.32 ;
    RECT 40.03 0.0 42.92 0.32 ;
    RECT 39.245 0.0 39.61 0.32 ;
    RECT 38.3 0.0 38.445 0.32 ;
    RECT 37.14 0.0 37.495 0.32 ;
    RECT 33.83 0.0 36.72 0.32 ;
    RECT 33.045 0.0 33.41 0.32 ;
    RECT 32.1 0.0 32.245 0.32 ;
    RECT 30.94 0.0 31.295 0.32 ;
    RECT 27.63 0.0 30.52 0.32 ;
    RECT 26.845 0.0 27.21 0.32 ;
    RECT 25.9 0.0 26.045 0.32 ;
    RECT 24.74 0.0 25.095 0.32 ;
    RECT 21.43 0.0 24.32 0.32 ;
    RECT 20.645 0.0 21.01 0.32 ;
    RECT 19.7 0.0 19.845 0.32 ;
    RECT 18.54 0.0 18.895 0.32 ;
    RECT 15.23 0.0 18.12 0.32 ;
    RECT 14.445 0.0 14.81 0.32 ;
    RECT 13.5 0.0 13.645 0.32 ;
    RECT 12.34 0.0 12.695 0.32 ;
    RECT 9.03 0.0 11.92 0.32 ;
    RECT 8.245 0.0 8.61 0.32 ;
    RECT 7.3 0.0 7.445 0.32 ;
    RECT 6.14 0.0 6.495 0.32 ;
    RECT 2.83 0.0 5.72 0.32 ;
    RECT 2.045 0.0 2.41 0.32 ;
    RECT 0.7 0.0 0.84 0.32 ;
    RECT 0.0 0.0 0.28 0.32 ;
    RECT 0.0 0.32 442.43 69.945 ;
    LAYER V2 ;
    RECT 0.0 0.0 442.43 69.945 ;
    LAYER M3 DESIGNRULEWIDTH 0.07 ;
    RECT 442.15 0.0 442.43 0.32 ;
    RECT 441.59 0.0 441.73 0.32 ;
    RECT 440.02 0.0 440.385 0.32 ;
    RECT 436.71 0.0 439.6 0.32 ;
    RECT 435.935 0.0 436.29 0.32 ;
    RECT 434.985 0.0 435.13 0.32 ;
    RECT 433.82 0.0 434.185 0.32 ;
    RECT 430.51 0.0 433.4 0.32 ;
    RECT 429.735 0.0 430.09 0.32 ;
    RECT 428.785 0.0 428.93 0.32 ;
    RECT 427.62 0.0 427.985 0.32 ;
    RECT 424.31 0.0 427.2 0.32 ;
    RECT 423.535 0.0 423.89 0.32 ;
    RECT 422.585 0.0 422.73 0.32 ;
    RECT 421.42 0.0 421.785 0.32 ;
    RECT 418.11 0.0 421.0 0.32 ;
    RECT 417.335 0.0 417.69 0.32 ;
    RECT 416.385 0.0 416.53 0.32 ;
    RECT 415.22 0.0 415.585 0.32 ;
    RECT 411.91 0.0 414.8 0.32 ;
    RECT 411.135 0.0 411.49 0.32 ;
    RECT 410.185 0.0 410.33 0.32 ;
    RECT 409.02 0.0 409.385 0.32 ;
    RECT 405.71 0.0 408.6 0.32 ;
    RECT 404.935 0.0 405.29 0.32 ;
    RECT 403.985 0.0 404.13 0.32 ;
    RECT 402.82 0.0 403.185 0.32 ;
    RECT 399.51 0.0 402.4 0.32 ;
    RECT 398.735 0.0 399.09 0.32 ;
    RECT 397.785 0.0 397.93 0.32 ;
    RECT 396.62 0.0 396.985 0.32 ;
    RECT 393.31 0.0 396.2 0.32 ;
    RECT 392.535 0.0 392.89 0.32 ;
    RECT 391.585 0.0 391.73 0.32 ;
    RECT 390.42 0.0 390.785 0.32 ;
    RECT 387.11 0.0 390.0 0.32 ;
    RECT 386.335 0.0 386.69 0.32 ;
    RECT 385.385 0.0 385.53 0.32 ;
    RECT 384.22 0.0 384.585 0.32 ;
    RECT 380.91 0.0 383.8 0.32 ;
    RECT 380.135 0.0 380.49 0.32 ;
    RECT 379.185 0.0 379.33 0.32 ;
    RECT 378.02 0.0 378.385 0.32 ;
    RECT 374.71 0.0 377.6 0.32 ;
    RECT 373.935 0.0 374.29 0.32 ;
    RECT 372.985 0.0 373.13 0.32 ;
    RECT 371.82 0.0 372.185 0.32 ;
    RECT 368.51 0.0 371.4 0.32 ;
    RECT 367.735 0.0 368.09 0.32 ;
    RECT 366.785 0.0 366.93 0.32 ;
    RECT 365.62 0.0 365.985 0.32 ;
    RECT 362.31 0.0 365.2 0.32 ;
    RECT 361.535 0.0 361.89 0.32 ;
    RECT 360.585 0.0 360.73 0.32 ;
    RECT 359.42 0.0 359.785 0.32 ;
    RECT 356.11 0.0 359.0 0.32 ;
    RECT 355.335 0.0 355.69 0.32 ;
    RECT 354.385 0.0 354.53 0.32 ;
    RECT 353.22 0.0 353.585 0.32 ;
    RECT 349.91 0.0 352.8 0.32 ;
    RECT 349.135 0.0 349.49 0.32 ;
    RECT 348.185 0.0 348.33 0.32 ;
    RECT 347.02 0.0 347.385 0.32 ;
    RECT 343.71 0.0 346.6 0.32 ;
    RECT 342.935 0.0 343.29 0.32 ;
    RECT 341.985 0.0 342.13 0.32 ;
    RECT 340.82 0.0 341.185 0.32 ;
    RECT 337.51 0.0 340.4 0.32 ;
    RECT 336.735 0.0 337.09 0.32 ;
    RECT 335.785 0.0 335.93 0.32 ;
    RECT 334.62 0.0 334.985 0.32 ;
    RECT 331.31 0.0 334.2 0.32 ;
    RECT 330.535 0.0 330.89 0.32 ;
    RECT 329.585 0.0 329.73 0.32 ;
    RECT 328.42 0.0 328.785 0.32 ;
    RECT 325.11 0.0 328.0 0.32 ;
    RECT 324.335 0.0 324.69 0.32 ;
    RECT 323.385 0.0 323.53 0.32 ;
    RECT 322.22 0.0 322.585 0.32 ;
    RECT 318.91 0.0 321.8 0.32 ;
    RECT 318.135 0.0 318.49 0.32 ;
    RECT 317.185 0.0 317.33 0.32 ;
    RECT 316.02 0.0 316.385 0.32 ;
    RECT 312.71 0.0 315.6 0.32 ;
    RECT 311.935 0.0 312.29 0.32 ;
    RECT 310.985 0.0 311.13 0.32 ;
    RECT 309.82 0.0 310.185 0.32 ;
    RECT 306.51 0.0 309.4 0.32 ;
    RECT 305.735 0.0 306.09 0.32 ;
    RECT 304.785 0.0 304.93 0.32 ;
    RECT 303.62 0.0 303.985 0.32 ;
    RECT 300.31 0.0 303.2 0.32 ;
    RECT 299.535 0.0 299.89 0.32 ;
    RECT 298.585 0.0 298.73 0.32 ;
    RECT 297.42 0.0 297.785 0.32 ;
    RECT 294.11 0.0 297.0 0.32 ;
    RECT 293.335 0.0 293.69 0.32 ;
    RECT 290.27 0.0 291.395 0.32 ;
    RECT 289.485 0.0 289.85 0.32 ;
    RECT 287.905 0.0 288.78 0.32 ;
    RECT 287.345 0.0 287.485 0.32 ;
    RECT 286.775 0.0 286.925 0.32 ;
    RECT 286.215 0.0 286.355 0.32 ;
    RECT 285.615 0.0 285.795 0.32 ;
    RECT 281.535 0.0 284.805 0.32 ;
    RECT 280.125 0.0 280.27 0.32 ;
    RECT 279.415 0.0 279.705 0.32 ;
    RECT 276.665 0.0 278.645 0.32 ;
    RECT 274.945 0.0 276.245 0.32 ;
    RECT 273.8 0.0 273.95 0.32 ;
    RECT 273.215 0.0 273.38 0.32 ;
    RECT 271.605 0.0 272.405 0.32 ;
    RECT 270.635 0.0 270.905 0.32 ;
    RECT 269.135 0.0 270.215 0.32 ;
    RECT 263.105 0.0 266.205 0.32 ;
    RECT 262.545 0.0 262.685 0.32 ;
    RECT 262.015 0.0 262.125 0.32 ;
    RECT 257.875 0.0 259.705 0.32 ;
    RECT 257.025 0.0 257.455 0.32 ;
    RECT 255.215 0.0 255.365 0.32 ;
    RECT 254.615 0.0 254.795 0.32 ;
    RECT 253.16 0.0 253.805 0.32 ;
    RECT 252.1 0.0 252.445 0.32 ;
    RECT 250.575 0.0 251.38 0.32 ;
    RECT 249.66 0.0 249.86 0.32 ;
    RECT 249.095 0.0 249.24 0.32 ;
    RECT 248.415 0.0 248.675 0.32 ;
    RECT 244.315 0.0 247.605 0.32 ;
    RECT 241.54 0.0 242.565 0.32 ;
    RECT 240.985 0.0 241.12 0.32 ;
    RECT 239.93 0.0 240.13 0.32 ;
    RECT 238.05 0.0 239.13 0.32 ;
    RECT 235.96 0.0 237.22 0.32 ;
    RECT 231.965 0.0 235.095 0.32 ;
    RECT 231.3 0.0 231.545 0.32 ;
    RECT 222.235 0.0 230.88 0.32 ;
    RECT 211.79 0.0 221.815 0.32 ;
    RECT 210.885 0.0 211.07 0.32 ;
    RECT 207.31 0.0 210.465 0.32 ;
    RECT 206.57 0.0 206.89 0.32 ;
    RECT 205.845 0.0 206.15 0.32 ;
    RECT 203.3 0.0 205.12 0.32 ;
    RECT 202.105 0.0 202.5 0.32 ;
    RECT 201.505 0.0 201.685 0.32 ;
    RECT 200.08 0.0 200.635 0.32 ;
    RECT 199.465 0.0 199.66 0.32 ;
    RECT 194.825 0.0 198.135 0.32 ;
    RECT 193.965 0.0 194.105 0.32 ;
    RECT 193.405 0.0 193.545 0.32 ;
    RECT 192.705 0.0 192.985 0.32 ;
    RECT 190.785 0.0 191.895 0.32 ;
    RECT 188.625 0.0 189.39 0.32 ;
    RECT 187.62 0.0 187.815 0.32 ;
    RECT 184.91 0.0 185.5 0.32 ;
    RECT 182.66 0.0 184.49 0.32 ;
    RECT 179.555 0.0 179.84 0.32 ;
    RECT 176.225 0.0 179.135 0.32 ;
    RECT 171.99 0.0 173.295 0.32 ;
    RECT 171.445 0.0 171.57 0.32 ;
    RECT 170.025 0.0 170.725 0.32 ;
    RECT 169.075 0.0 169.215 0.32 ;
    RECT 168.505 0.0 168.655 0.32 ;
    RECT 167.255 0.0 167.445 0.32 ;
    RECT 166.215 0.0 166.835 0.32 ;
    RECT 163.775 0.0 165.795 0.32 ;
    RECT 162.895 0.0 163.045 0.32 ;
    RECT 162.305 0.0 162.475 0.32 ;
    RECT 161.705 0.0 161.885 0.32 ;
    RECT 157.625 0.0 160.895 0.32 ;
    RECT 156.275 0.0 156.435 0.32 ;
    RECT 155.34 0.0 155.855 0.32 ;
    RECT 153.795 0.0 154.92 0.32 ;
    RECT 152.65 0.0 153.0 0.32 ;
    RECT 151.72 0.0 152.23 0.32 ;
    RECT 151.035 0.0 151.3 0.32 ;
    RECT 149.9 0.0 150.035 0.32 ;
    RECT 148.74 0.0 149.095 0.32 ;
    RECT 145.43 0.0 148.32 0.32 ;
    RECT 144.645 0.0 145.01 0.32 ;
    RECT 143.7 0.0 143.845 0.32 ;
    RECT 142.54 0.0 142.895 0.32 ;
    RECT 139.23 0.0 142.12 0.32 ;
    RECT 138.445 0.0 138.81 0.32 ;
    RECT 137.5 0.0 137.645 0.32 ;
    RECT 136.34 0.0 136.695 0.32 ;
    RECT 133.03 0.0 135.92 0.32 ;
    RECT 132.245 0.0 132.61 0.32 ;
    RECT 131.3 0.0 131.445 0.32 ;
    RECT 130.14 0.0 130.495 0.32 ;
    RECT 126.83 0.0 129.72 0.32 ;
    RECT 126.045 0.0 126.41 0.32 ;
    RECT 125.1 0.0 125.245 0.32 ;
    RECT 123.94 0.0 124.295 0.32 ;
    RECT 120.63 0.0 123.52 0.32 ;
    RECT 119.845 0.0 120.21 0.32 ;
    RECT 118.9 0.0 119.045 0.32 ;
    RECT 117.74 0.0 118.095 0.32 ;
    RECT 114.43 0.0 117.32 0.32 ;
    RECT 113.645 0.0 114.01 0.32 ;
    RECT 112.7 0.0 112.845 0.32 ;
    RECT 111.54 0.0 111.895 0.32 ;
    RECT 108.23 0.0 111.12 0.32 ;
    RECT 107.445 0.0 107.81 0.32 ;
    RECT 106.5 0.0 106.645 0.32 ;
    RECT 105.34 0.0 105.695 0.32 ;
    RECT 102.03 0.0 104.92 0.32 ;
    RECT 101.245 0.0 101.61 0.32 ;
    RECT 100.3 0.0 100.445 0.32 ;
    RECT 99.14 0.0 99.495 0.32 ;
    RECT 95.83 0.0 98.72 0.32 ;
    RECT 95.045 0.0 95.41 0.32 ;
    RECT 94.1 0.0 94.245 0.32 ;
    RECT 92.94 0.0 93.295 0.32 ;
    RECT 89.63 0.0 92.52 0.32 ;
    RECT 88.845 0.0 89.21 0.32 ;
    RECT 87.9 0.0 88.045 0.32 ;
    RECT 86.74 0.0 87.095 0.32 ;
    RECT 83.43 0.0 86.32 0.32 ;
    RECT 82.645 0.0 83.01 0.32 ;
    RECT 81.7 0.0 81.845 0.32 ;
    RECT 80.54 0.0 80.895 0.32 ;
    RECT 77.23 0.0 80.12 0.32 ;
    RECT 76.445 0.0 76.81 0.32 ;
    RECT 75.5 0.0 75.645 0.32 ;
    RECT 74.34 0.0 74.695 0.32 ;
    RECT 71.03 0.0 73.92 0.32 ;
    RECT 70.245 0.0 70.61 0.32 ;
    RECT 69.3 0.0 69.445 0.32 ;
    RECT 68.14 0.0 68.495 0.32 ;
    RECT 64.83 0.0 67.72 0.32 ;
    RECT 64.045 0.0 64.41 0.32 ;
    RECT 63.1 0.0 63.245 0.32 ;
    RECT 61.94 0.0 62.295 0.32 ;
    RECT 58.63 0.0 61.52 0.32 ;
    RECT 57.845 0.0 58.21 0.32 ;
    RECT 56.9 0.0 57.045 0.32 ;
    RECT 55.74 0.0 56.095 0.32 ;
    RECT 52.43 0.0 55.32 0.32 ;
    RECT 51.645 0.0 52.01 0.32 ;
    RECT 50.7 0.0 50.845 0.32 ;
    RECT 49.54 0.0 49.895 0.32 ;
    RECT 46.23 0.0 49.12 0.32 ;
    RECT 45.445 0.0 45.81 0.32 ;
    RECT 44.5 0.0 44.645 0.32 ;
    RECT 43.34 0.0 43.695 0.32 ;
    RECT 40.03 0.0 42.92 0.32 ;
    RECT 39.245 0.0 39.61 0.32 ;
    RECT 38.3 0.0 38.445 0.32 ;
    RECT 37.14 0.0 37.495 0.32 ;
    RECT 33.83 0.0 36.72 0.32 ;
    RECT 33.045 0.0 33.41 0.32 ;
    RECT 32.1 0.0 32.245 0.32 ;
    RECT 30.94 0.0 31.295 0.32 ;
    RECT 27.63 0.0 30.52 0.32 ;
    RECT 26.845 0.0 27.21 0.32 ;
    RECT 25.9 0.0 26.045 0.32 ;
    RECT 24.74 0.0 25.095 0.32 ;
    RECT 21.43 0.0 24.32 0.32 ;
    RECT 20.645 0.0 21.01 0.32 ;
    RECT 19.7 0.0 19.845 0.32 ;
    RECT 18.54 0.0 18.895 0.32 ;
    RECT 15.23 0.0 18.12 0.32 ;
    RECT 14.445 0.0 14.81 0.32 ;
    RECT 13.5 0.0 13.645 0.32 ;
    RECT 12.34 0.0 12.695 0.32 ;
    RECT 9.03 0.0 11.92 0.32 ;
    RECT 8.245 0.0 8.61 0.32 ;
    RECT 7.3 0.0 7.445 0.32 ;
    RECT 6.14 0.0 6.495 0.32 ;
    RECT 2.83 0.0 5.72 0.32 ;
    RECT 2.045 0.0 2.41 0.32 ;
    RECT 0.7 0.0 0.84 0.32 ;
    RECT 0.0 0.0 0.28 0.32 ;
    RECT 0.0 0.32 442.43 69.945 ;
    LAYER V3 ;
    RECT 0.0 0.0 442.43 69.945 ;
    LAYER M4 DESIGNRULEWIDTH 0.07 ;
    RECT 441.445 0.0 442.43 0.32 ;
    RECT 440.875 0.0 441.095 0.32 ;
    RECT 439.895 0.0 440.525 0.32 ;
    RECT 438.345 0.0 439.545 0.32 ;
    RECT 437.765 0.0 437.995 0.32 ;
    RECT 436.795 0.0 437.415 0.32 ;
    RECT 435.815 0.0 436.445 0.32 ;
    RECT 435.245 0.0 435.465 0.32 ;
    RECT 434.675 0.0 434.895 0.32 ;
    RECT 433.695 0.0 434.325 0.32 ;
    RECT 432.145 0.0 433.345 0.32 ;
    RECT 431.565 0.0 431.795 0.32 ;
    RECT 430.595 0.0 431.215 0.32 ;
    RECT 429.615 0.0 430.245 0.32 ;
    RECT 429.045 0.0 429.265 0.32 ;
    RECT 428.475 0.0 428.695 0.32 ;
    RECT 427.495 0.0 428.125 0.32 ;
    RECT 425.945 0.0 427.145 0.32 ;
    RECT 425.365 0.0 425.595 0.32 ;
    RECT 424.395 0.0 425.015 0.32 ;
    RECT 423.415 0.0 424.045 0.32 ;
    RECT 422.845 0.0 423.065 0.32 ;
    RECT 422.275 0.0 422.495 0.32 ;
    RECT 421.295 0.0 421.925 0.32 ;
    RECT 419.745 0.0 420.945 0.32 ;
    RECT 419.165 0.0 419.395 0.32 ;
    RECT 418.195 0.0 418.815 0.32 ;
    RECT 417.215 0.0 417.845 0.32 ;
    RECT 416.645 0.0 416.865 0.32 ;
    RECT 416.075 0.0 416.295 0.32 ;
    RECT 415.095 0.0 415.725 0.32 ;
    RECT 413.545 0.0 414.745 0.32 ;
    RECT 412.965 0.0 413.195 0.32 ;
    RECT 411.995 0.0 412.615 0.32 ;
    RECT 411.015 0.0 411.645 0.32 ;
    RECT 410.445 0.0 410.665 0.32 ;
    RECT 409.875 0.0 410.095 0.32 ;
    RECT 408.895 0.0 409.525 0.32 ;
    RECT 407.345 0.0 408.545 0.32 ;
    RECT 406.765 0.0 406.995 0.32 ;
    RECT 405.795 0.0 406.415 0.32 ;
    RECT 404.815 0.0 405.445 0.32 ;
    RECT 404.245 0.0 404.465 0.32 ;
    RECT 403.675 0.0 403.895 0.32 ;
    RECT 402.695 0.0 403.325 0.32 ;
    RECT 401.145 0.0 402.345 0.32 ;
    RECT 400.565 0.0 400.795 0.32 ;
    RECT 399.595 0.0 400.215 0.32 ;
    RECT 398.615 0.0 399.245 0.32 ;
    RECT 398.045 0.0 398.265 0.32 ;
    RECT 397.475 0.0 397.695 0.32 ;
    RECT 396.495 0.0 397.125 0.32 ;
    RECT 394.945 0.0 396.145 0.32 ;
    RECT 394.365 0.0 394.595 0.32 ;
    RECT 393.395 0.0 394.015 0.32 ;
    RECT 392.415 0.0 393.045 0.32 ;
    RECT 391.845 0.0 392.065 0.32 ;
    RECT 391.275 0.0 391.495 0.32 ;
    RECT 390.295 0.0 390.925 0.32 ;
    RECT 388.745 0.0 389.945 0.32 ;
    RECT 388.165 0.0 388.395 0.32 ;
    RECT 387.195 0.0 387.815 0.32 ;
    RECT 386.215 0.0 386.845 0.32 ;
    RECT 385.645 0.0 385.865 0.32 ;
    RECT 385.075 0.0 385.295 0.32 ;
    RECT 384.095 0.0 384.725 0.32 ;
    RECT 382.545 0.0 383.745 0.32 ;
    RECT 381.965 0.0 382.195 0.32 ;
    RECT 380.995 0.0 381.615 0.32 ;
    RECT 380.015 0.0 380.645 0.32 ;
    RECT 379.445 0.0 379.665 0.32 ;
    RECT 378.875 0.0 379.095 0.32 ;
    RECT 377.895 0.0 378.525 0.32 ;
    RECT 376.345 0.0 377.545 0.32 ;
    RECT 375.765 0.0 375.995 0.32 ;
    RECT 374.795 0.0 375.415 0.32 ;
    RECT 373.815 0.0 374.445 0.32 ;
    RECT 373.245 0.0 373.465 0.32 ;
    RECT 372.675 0.0 372.895 0.32 ;
    RECT 371.695 0.0 372.325 0.32 ;
    RECT 370.145 0.0 371.345 0.32 ;
    RECT 369.565 0.0 369.795 0.32 ;
    RECT 368.595 0.0 369.215 0.32 ;
    RECT 367.615 0.0 368.245 0.32 ;
    RECT 367.045 0.0 367.265 0.32 ;
    RECT 366.475 0.0 366.695 0.32 ;
    RECT 365.495 0.0 366.125 0.32 ;
    RECT 363.945 0.0 365.145 0.32 ;
    RECT 363.365 0.0 363.595 0.32 ;
    RECT 362.395 0.0 363.015 0.32 ;
    RECT 361.415 0.0 362.045 0.32 ;
    RECT 360.845 0.0 361.065 0.32 ;
    RECT 360.275 0.0 360.495 0.32 ;
    RECT 359.295 0.0 359.925 0.32 ;
    RECT 357.745 0.0 358.945 0.32 ;
    RECT 357.165 0.0 357.395 0.32 ;
    RECT 356.195 0.0 356.815 0.32 ;
    RECT 355.215 0.0 355.845 0.32 ;
    RECT 354.645 0.0 354.865 0.32 ;
    RECT 354.075 0.0 354.295 0.32 ;
    RECT 353.095 0.0 353.725 0.32 ;
    RECT 351.545 0.0 352.745 0.32 ;
    RECT 350.965 0.0 351.195 0.32 ;
    RECT 349.995 0.0 350.615 0.32 ;
    RECT 349.015 0.0 349.645 0.32 ;
    RECT 348.445 0.0 348.665 0.32 ;
    RECT 347.875 0.0 348.095 0.32 ;
    RECT 346.895 0.0 347.525 0.32 ;
    RECT 345.345 0.0 346.545 0.32 ;
    RECT 344.765 0.0 344.995 0.32 ;
    RECT 343.795 0.0 344.415 0.32 ;
    RECT 342.815 0.0 343.445 0.32 ;
    RECT 342.245 0.0 342.465 0.32 ;
    RECT 341.675 0.0 341.895 0.32 ;
    RECT 340.695 0.0 341.325 0.32 ;
    RECT 339.145 0.0 340.345 0.32 ;
    RECT 338.565 0.0 338.795 0.32 ;
    RECT 337.595 0.0 338.215 0.32 ;
    RECT 336.615 0.0 337.245 0.32 ;
    RECT 336.045 0.0 336.265 0.32 ;
    RECT 335.475 0.0 335.695 0.32 ;
    RECT 334.495 0.0 335.125 0.32 ;
    RECT 332.945 0.0 334.145 0.32 ;
    RECT 332.365 0.0 332.595 0.32 ;
    RECT 331.395 0.0 332.015 0.32 ;
    RECT 330.415 0.0 331.045 0.32 ;
    RECT 329.845 0.0 330.065 0.32 ;
    RECT 329.275 0.0 329.495 0.32 ;
    RECT 328.295 0.0 328.925 0.32 ;
    RECT 326.745 0.0 327.945 0.32 ;
    RECT 326.165 0.0 326.395 0.32 ;
    RECT 325.195 0.0 325.815 0.32 ;
    RECT 324.215 0.0 324.845 0.32 ;
    RECT 323.645 0.0 323.865 0.32 ;
    RECT 323.075 0.0 323.295 0.32 ;
    RECT 322.095 0.0 322.725 0.32 ;
    RECT 320.545 0.0 321.745 0.32 ;
    RECT 319.965 0.0 320.195 0.32 ;
    RECT 318.995 0.0 319.615 0.32 ;
    RECT 318.015 0.0 318.645 0.32 ;
    RECT 317.445 0.0 317.665 0.32 ;
    RECT 316.875 0.0 317.095 0.32 ;
    RECT 315.895 0.0 316.525 0.32 ;
    RECT 314.345 0.0 315.545 0.32 ;
    RECT 313.765 0.0 313.995 0.32 ;
    RECT 312.795 0.0 313.415 0.32 ;
    RECT 311.815 0.0 312.445 0.32 ;
    RECT 311.245 0.0 311.465 0.32 ;
    RECT 310.675 0.0 310.895 0.32 ;
    RECT 309.695 0.0 310.325 0.32 ;
    RECT 308.145 0.0 309.345 0.32 ;
    RECT 307.565 0.0 307.795 0.32 ;
    RECT 306.595 0.0 307.215 0.32 ;
    RECT 305.615 0.0 306.245 0.32 ;
    RECT 305.045 0.0 305.265 0.32 ;
    RECT 304.475 0.0 304.695 0.32 ;
    RECT 303.495 0.0 304.125 0.32 ;
    RECT 301.945 0.0 303.145 0.32 ;
    RECT 301.365 0.0 301.595 0.32 ;
    RECT 300.395 0.0 301.015 0.32 ;
    RECT 299.415 0.0 300.045 0.32 ;
    RECT 298.845 0.0 299.065 0.32 ;
    RECT 298.275 0.0 298.495 0.32 ;
    RECT 297.295 0.0 297.925 0.32 ;
    RECT 295.745 0.0 296.945 0.32 ;
    RECT 295.165 0.0 295.395 0.32 ;
    RECT 294.195 0.0 294.815 0.32 ;
    RECT 293.215 0.0 293.845 0.32 ;
    RECT 292.645 0.0 292.865 0.32 ;
    RECT 292.075 0.0 292.295 0.32 ;
    RECT 291.095 0.0 291.395 0.32 ;
    RECT 289.545 0.0 290.745 0.32 ;
    RECT 288.965 0.0 289.195 0.32 ;
    RECT 287.995 0.0 288.615 0.32 ;
    RECT 287.345 0.0 287.645 0.32 ;
    RECT 286.445 0.0 286.665 0.32 ;
    RECT 285.875 0.0 286.095 0.32 ;
    RECT 283.345 0.0 284.545 0.32 ;
    RECT 282.765 0.0 282.995 0.32 ;
    RECT 281.795 0.0 282.415 0.32 ;
    RECT 280.245 0.0 280.465 0.32 ;
    RECT 279.675 0.0 279.895 0.32 ;
    RECT 278.695 0.0 278.995 0.32 ;
    RECT 277.145 0.0 278.345 0.32 ;
    RECT 276.565 0.0 276.795 0.32 ;
    RECT 275.595 0.0 276.215 0.32 ;
    RECT 274.945 0.0 275.245 0.32 ;
    RECT 274.045 0.0 274.265 0.32 ;
    RECT 273.475 0.0 273.695 0.32 ;
    RECT 270.945 0.0 272.145 0.32 ;
    RECT 270.365 0.0 270.595 0.32 ;
    RECT 269.395 0.0 270.015 0.32 ;
    RECT 267.845 0.0 268.065 0.32 ;
    RECT 267.275 0.0 267.495 0.32 ;
    RECT 264.745 0.0 265.945 0.32 ;
    RECT 264.165 0.0 264.395 0.32 ;
    RECT 263.195 0.0 263.815 0.32 ;
    RECT 262.545 0.0 262.845 0.32 ;
    RECT 261.645 0.0 261.865 0.32 ;
    RECT 261.075 0.0 261.295 0.32 ;
    RECT 258.545 0.0 259.745 0.32 ;
    RECT 257.965 0.0 258.195 0.32 ;
    RECT 256.995 0.0 257.615 0.32 ;
    RECT 255.445 0.0 255.665 0.32 ;
    RECT 254.875 0.0 255.095 0.32 ;
    RECT 252.345 0.0 253.545 0.32 ;
    RECT 251.765 0.0 251.995 0.32 ;
    RECT 250.795 0.0 251.415 0.32 ;
    RECT 250.28 0.0 250.445 0.32 ;
    RECT 249.245 0.0 249.465 0.32 ;
    RECT 248.675 0.0 248.895 0.32 ;
    RECT 246.145 0.0 247.345 0.32 ;
    RECT 245.565 0.0 245.795 0.32 ;
    RECT 244.595 0.0 245.215 0.32 ;
    RECT 243.945 0.0 244.245 0.32 ;
    RECT 243.045 0.0 243.265 0.32 ;
    RECT 241.305 0.0 242.695 0.32 ;
    RECT 240.515 0.0 240.955 0.32 ;
    RECT 239.515 0.0 240.165 0.32 ;
    RECT 235.96 0.0 236.82 0.32 ;
    RECT 235.4 0.0 235.48 0.32 ;
    RECT 233.84 0.0 234.27 0.32 ;
    RECT 232.705 0.0 233.49 0.32 ;
    RECT 231.965 0.0 232.225 0.32 ;
    RECT 231.44 0.0 231.545 0.32 ;
    RECT 230.675 0.0 230.98 0.32 ;
    RECT 229.505 0.0 229.935 0.32 ;
    RECT 227.565 0.0 227.995 0.32 ;
    RECT 226.915 0.0 227.215 0.32 ;
    RECT 225.32 0.0 225.79 0.32 ;
    RECT 224.52 0.0 224.97 0.32 ;
    RECT 223.95 0.0 224.17 0.32 ;
    RECT 222.29 0.0 223.49 0.32 ;
    RECT 221.78 0.0 221.94 0.32 ;
    RECT 221.0 0.0 221.43 0.32 ;
    RECT 220.49 0.0 220.65 0.32 ;
    RECT 218.94 0.0 220.14 0.32 ;
    RECT 218.26 0.0 218.48 0.32 ;
    RECT 217.46 0.0 217.91 0.32 ;
    RECT 216.64 0.0 217.11 0.32 ;
    RECT 215.215 0.0 215.515 0.32 ;
    RECT 214.435 0.0 214.865 0.32 ;
    RECT 212.495 0.0 212.925 0.32 ;
    RECT 210.885 0.0 210.99 0.32 ;
    RECT 210.205 0.0 210.465 0.32 ;
    RECT 208.94 0.0 209.725 0.32 ;
    RECT 208.16 0.0 208.59 0.32 ;
    RECT 206.95 0.0 207.03 0.32 ;
    RECT 205.61 0.0 206.47 0.32 ;
    RECT 202.265 0.0 202.915 0.32 ;
    RECT 201.475 0.0 201.915 0.32 ;
    RECT 199.735 0.0 201.125 0.32 ;
    RECT 199.165 0.0 199.385 0.32 ;
    RECT 198.185 0.0 198.485 0.32 ;
    RECT 197.215 0.0 197.835 0.32 ;
    RECT 196.635 0.0 196.865 0.32 ;
    RECT 195.085 0.0 196.285 0.32 ;
    RECT 193.535 0.0 193.755 0.32 ;
    RECT 192.965 0.0 193.185 0.32 ;
    RECT 191.015 0.0 191.635 0.32 ;
    RECT 190.435 0.0 190.665 0.32 ;
    RECT 188.885 0.0 190.085 0.32 ;
    RECT 187.335 0.0 187.555 0.32 ;
    RECT 186.765 0.0 186.985 0.32 ;
    RECT 184.815 0.0 185.435 0.32 ;
    RECT 184.235 0.0 184.465 0.32 ;
    RECT 182.685 0.0 183.885 0.32 ;
    RECT 181.135 0.0 181.355 0.32 ;
    RECT 180.565 0.0 180.785 0.32 ;
    RECT 179.585 0.0 179.84 0.32 ;
    RECT 178.615 0.0 179.235 0.32 ;
    RECT 178.035 0.0 178.265 0.32 ;
    RECT 176.485 0.0 177.685 0.32 ;
    RECT 174.935 0.0 175.155 0.32 ;
    RECT 174.365 0.0 174.585 0.32 ;
    RECT 172.415 0.0 173.035 0.32 ;
    RECT 171.835 0.0 172.065 0.32 ;
    RECT 170.285 0.0 171.485 0.32 ;
    RECT 168.735 0.0 168.955 0.32 ;
    RECT 168.165 0.0 168.385 0.32 ;
    RECT 167.185 0.0 167.445 0.32 ;
    RECT 166.215 0.0 166.835 0.32 ;
    RECT 165.635 0.0 165.865 0.32 ;
    RECT 164.085 0.0 165.285 0.32 ;
    RECT 163.465 0.0 163.735 0.32 ;
    RECT 162.535 0.0 162.755 0.32 ;
    RECT 161.965 0.0 162.185 0.32 ;
    RECT 160.015 0.0 160.635 0.32 ;
    RECT 159.435 0.0 159.665 0.32 ;
    RECT 157.885 0.0 159.085 0.32 ;
    RECT 156.335 0.0 156.555 0.32 ;
    RECT 155.765 0.0 155.985 0.32 ;
    RECT 155.34 0.0 155.415 0.32 ;
    RECT 154.785 0.0 154.92 0.32 ;
    RECT 153.815 0.0 154.435 0.32 ;
    RECT 153.235 0.0 153.465 0.32 ;
    RECT 151.685 0.0 152.885 0.32 ;
    RECT 151.035 0.0 151.335 0.32 ;
    RECT 150.135 0.0 150.355 0.32 ;
    RECT 149.565 0.0 149.785 0.32 ;
    RECT 148.585 0.0 149.215 0.32 ;
    RECT 147.615 0.0 148.235 0.32 ;
    RECT 147.035 0.0 147.265 0.32 ;
    RECT 145.485 0.0 146.685 0.32 ;
    RECT 144.505 0.0 145.135 0.32 ;
    RECT 143.935 0.0 144.155 0.32 ;
    RECT 143.365 0.0 143.585 0.32 ;
    RECT 142.385 0.0 143.015 0.32 ;
    RECT 141.415 0.0 142.035 0.32 ;
    RECT 140.835 0.0 141.065 0.32 ;
    RECT 139.285 0.0 140.485 0.32 ;
    RECT 138.305 0.0 138.935 0.32 ;
    RECT 137.735 0.0 137.955 0.32 ;
    RECT 137.165 0.0 137.385 0.32 ;
    RECT 136.185 0.0 136.815 0.32 ;
    RECT 135.215 0.0 135.835 0.32 ;
    RECT 134.635 0.0 134.865 0.32 ;
    RECT 133.085 0.0 134.285 0.32 ;
    RECT 132.105 0.0 132.735 0.32 ;
    RECT 131.535 0.0 131.755 0.32 ;
    RECT 130.965 0.0 131.185 0.32 ;
    RECT 129.985 0.0 130.615 0.32 ;
    RECT 129.015 0.0 129.635 0.32 ;
    RECT 128.435 0.0 128.665 0.32 ;
    RECT 126.885 0.0 128.085 0.32 ;
    RECT 125.905 0.0 126.535 0.32 ;
    RECT 125.335 0.0 125.555 0.32 ;
    RECT 124.765 0.0 124.985 0.32 ;
    RECT 123.785 0.0 124.415 0.32 ;
    RECT 122.815 0.0 123.435 0.32 ;
    RECT 122.235 0.0 122.465 0.32 ;
    RECT 120.685 0.0 121.885 0.32 ;
    RECT 119.705 0.0 120.335 0.32 ;
    RECT 119.135 0.0 119.355 0.32 ;
    RECT 118.565 0.0 118.785 0.32 ;
    RECT 117.585 0.0 118.215 0.32 ;
    RECT 116.615 0.0 117.235 0.32 ;
    RECT 116.035 0.0 116.265 0.32 ;
    RECT 114.485 0.0 115.685 0.32 ;
    RECT 113.505 0.0 114.135 0.32 ;
    RECT 112.935 0.0 113.155 0.32 ;
    RECT 112.365 0.0 112.585 0.32 ;
    RECT 111.385 0.0 112.015 0.32 ;
    RECT 110.415 0.0 111.035 0.32 ;
    RECT 109.835 0.0 110.065 0.32 ;
    RECT 108.285 0.0 109.485 0.32 ;
    RECT 107.305 0.0 107.935 0.32 ;
    RECT 106.735 0.0 106.955 0.32 ;
    RECT 106.165 0.0 106.385 0.32 ;
    RECT 105.185 0.0 105.815 0.32 ;
    RECT 104.215 0.0 104.835 0.32 ;
    RECT 103.635 0.0 103.865 0.32 ;
    RECT 102.085 0.0 103.285 0.32 ;
    RECT 101.105 0.0 101.735 0.32 ;
    RECT 100.535 0.0 100.755 0.32 ;
    RECT 99.965 0.0 100.185 0.32 ;
    RECT 98.985 0.0 99.615 0.32 ;
    RECT 98.015 0.0 98.635 0.32 ;
    RECT 97.435 0.0 97.665 0.32 ;
    RECT 95.885 0.0 97.085 0.32 ;
    RECT 94.905 0.0 95.535 0.32 ;
    RECT 94.335 0.0 94.555 0.32 ;
    RECT 93.765 0.0 93.985 0.32 ;
    RECT 92.785 0.0 93.415 0.32 ;
    RECT 91.815 0.0 92.435 0.32 ;
    RECT 91.235 0.0 91.465 0.32 ;
    RECT 89.685 0.0 90.885 0.32 ;
    RECT 88.705 0.0 89.335 0.32 ;
    RECT 88.135 0.0 88.355 0.32 ;
    RECT 87.565 0.0 87.785 0.32 ;
    RECT 86.585 0.0 87.215 0.32 ;
    RECT 85.615 0.0 86.235 0.32 ;
    RECT 85.035 0.0 85.265 0.32 ;
    RECT 83.485 0.0 84.685 0.32 ;
    RECT 82.505 0.0 83.135 0.32 ;
    RECT 81.935 0.0 82.155 0.32 ;
    RECT 81.365 0.0 81.585 0.32 ;
    RECT 80.385 0.0 81.015 0.32 ;
    RECT 79.415 0.0 80.035 0.32 ;
    RECT 78.835 0.0 79.065 0.32 ;
    RECT 77.285 0.0 78.485 0.32 ;
    RECT 76.305 0.0 76.935 0.32 ;
    RECT 75.735 0.0 75.955 0.32 ;
    RECT 75.165 0.0 75.385 0.32 ;
    RECT 74.185 0.0 74.815 0.32 ;
    RECT 73.215 0.0 73.835 0.32 ;
    RECT 72.635 0.0 72.865 0.32 ;
    RECT 71.085 0.0 72.285 0.32 ;
    RECT 70.105 0.0 70.735 0.32 ;
    RECT 69.535 0.0 69.755 0.32 ;
    RECT 68.965 0.0 69.185 0.32 ;
    RECT 67.985 0.0 68.615 0.32 ;
    RECT 67.015 0.0 67.635 0.32 ;
    RECT 66.435 0.0 66.665 0.32 ;
    RECT 64.885 0.0 66.085 0.32 ;
    RECT 63.905 0.0 64.535 0.32 ;
    RECT 63.335 0.0 63.555 0.32 ;
    RECT 62.765 0.0 62.985 0.32 ;
    RECT 61.785 0.0 62.415 0.32 ;
    RECT 60.815 0.0 61.435 0.32 ;
    RECT 60.235 0.0 60.465 0.32 ;
    RECT 58.685 0.0 59.885 0.32 ;
    RECT 57.705 0.0 58.335 0.32 ;
    RECT 57.135 0.0 57.355 0.32 ;
    RECT 56.565 0.0 56.785 0.32 ;
    RECT 55.585 0.0 56.215 0.32 ;
    RECT 54.615 0.0 55.235 0.32 ;
    RECT 54.035 0.0 54.265 0.32 ;
    RECT 52.485 0.0 53.685 0.32 ;
    RECT 51.505 0.0 52.135 0.32 ;
    RECT 50.935 0.0 51.155 0.32 ;
    RECT 50.365 0.0 50.585 0.32 ;
    RECT 49.385 0.0 50.015 0.32 ;
    RECT 48.415 0.0 49.035 0.32 ;
    RECT 47.835 0.0 48.065 0.32 ;
    RECT 46.285 0.0 47.485 0.32 ;
    RECT 45.305 0.0 45.935 0.32 ;
    RECT 44.735 0.0 44.955 0.32 ;
    RECT 44.165 0.0 44.385 0.32 ;
    RECT 43.185 0.0 43.815 0.32 ;
    RECT 42.215 0.0 42.835 0.32 ;
    RECT 41.635 0.0 41.865 0.32 ;
    RECT 40.085 0.0 41.285 0.32 ;
    RECT 39.105 0.0 39.735 0.32 ;
    RECT 38.535 0.0 38.755 0.32 ;
    RECT 37.965 0.0 38.185 0.32 ;
    RECT 36.985 0.0 37.615 0.32 ;
    RECT 36.015 0.0 36.635 0.32 ;
    RECT 35.435 0.0 35.665 0.32 ;
    RECT 33.885 0.0 35.085 0.32 ;
    RECT 32.905 0.0 33.535 0.32 ;
    RECT 32.335 0.0 32.555 0.32 ;
    RECT 31.765 0.0 31.985 0.32 ;
    RECT 30.785 0.0 31.415 0.32 ;
    RECT 29.815 0.0 30.435 0.32 ;
    RECT 29.235 0.0 29.465 0.32 ;
    RECT 27.685 0.0 28.885 0.32 ;
    RECT 26.705 0.0 27.335 0.32 ;
    RECT 26.135 0.0 26.355 0.32 ;
    RECT 25.565 0.0 25.785 0.32 ;
    RECT 24.585 0.0 25.215 0.32 ;
    RECT 23.615 0.0 24.235 0.32 ;
    RECT 23.035 0.0 23.265 0.32 ;
    RECT 21.485 0.0 22.685 0.32 ;
    RECT 20.505 0.0 21.135 0.32 ;
    RECT 19.935 0.0 20.155 0.32 ;
    RECT 19.365 0.0 19.585 0.32 ;
    RECT 18.385 0.0 19.015 0.32 ;
    RECT 17.415 0.0 18.035 0.32 ;
    RECT 16.835 0.0 17.065 0.32 ;
    RECT 15.285 0.0 16.485 0.32 ;
    RECT 14.305 0.0 14.935 0.32 ;
    RECT 13.735 0.0 13.955 0.32 ;
    RECT 13.165 0.0 13.385 0.32 ;
    RECT 12.185 0.0 12.815 0.32 ;
    RECT 11.215 0.0 11.835 0.32 ;
    RECT 10.635 0.0 10.865 0.32 ;
    RECT 9.085 0.0 10.285 0.32 ;
    RECT 8.105 0.0 8.735 0.32 ;
    RECT 7.535 0.0 7.755 0.32 ;
    RECT 6.965 0.0 7.185 0.32 ;
    RECT 5.985 0.0 6.615 0.32 ;
    RECT 5.015 0.0 5.635 0.32 ;
    RECT 4.435 0.0 4.665 0.32 ;
    RECT 2.885 0.0 4.085 0.32 ;
    RECT 1.905 0.0 2.535 0.32 ;
    RECT 1.335 0.0 1.555 0.32 ;
    RECT 0.0 0.0 0.985 0.32 ;
    RECT 441.445 0.32 442.43 69.945 ;
    RECT 440.875 0.32 441.095 69.945 ;
    RECT 439.895 0.32 440.525 69.945 ;
    RECT 438.345 0.32 439.545 69.945 ;
    RECT 437.765 0.32 437.995 69.945 ;
    RECT 436.795 0.32 437.415 69.945 ;
    RECT 435.815 0.32 436.445 69.945 ;
    RECT 435.245 0.32 435.465 69.945 ;
    RECT 434.675 0.32 434.895 69.945 ;
    RECT 433.695 0.32 434.325 69.945 ;
    RECT 432.145 0.32 433.345 69.945 ;
    RECT 431.565 0.32 431.795 69.945 ;
    RECT 430.595 0.32 431.215 69.945 ;
    RECT 429.615 0.32 430.245 69.945 ;
    RECT 429.045 0.32 429.265 69.945 ;
    RECT 428.475 0.32 428.695 69.945 ;
    RECT 427.495 0.32 428.125 69.945 ;
    RECT 425.945 0.32 427.145 69.945 ;
    RECT 425.365 0.32 425.595 69.945 ;
    RECT 424.395 0.32 425.015 69.945 ;
    RECT 423.415 0.32 424.045 69.945 ;
    RECT 422.845 0.32 423.065 69.945 ;
    RECT 422.275 0.32 422.495 69.945 ;
    RECT 421.295 0.32 421.925 69.945 ;
    RECT 419.745 0.32 420.945 69.945 ;
    RECT 419.165 0.32 419.395 69.945 ;
    RECT 418.195 0.32 418.815 69.945 ;
    RECT 417.215 0.32 417.845 69.945 ;
    RECT 416.645 0.32 416.865 69.945 ;
    RECT 416.075 0.32 416.295 69.945 ;
    RECT 415.095 0.32 415.725 69.945 ;
    RECT 413.545 0.32 414.745 69.945 ;
    RECT 412.965 0.32 413.195 69.945 ;
    RECT 411.995 0.32 412.615 69.945 ;
    RECT 411.015 0.32 411.645 69.945 ;
    RECT 410.445 0.32 410.665 69.945 ;
    RECT 409.875 0.32 410.095 69.945 ;
    RECT 408.895 0.32 409.525 69.945 ;
    RECT 407.345 0.32 408.545 69.945 ;
    RECT 406.765 0.32 406.995 69.945 ;
    RECT 405.795 0.32 406.415 69.945 ;
    RECT 404.815 0.32 405.445 69.945 ;
    RECT 404.245 0.32 404.465 69.945 ;
    RECT 403.675 0.32 403.895 69.945 ;
    RECT 402.695 0.32 403.325 69.945 ;
    RECT 401.145 0.32 402.345 69.945 ;
    RECT 400.565 0.32 400.795 69.945 ;
    RECT 399.595 0.32 400.215 69.945 ;
    RECT 398.615 0.32 399.245 69.945 ;
    RECT 398.045 0.32 398.265 69.945 ;
    RECT 397.475 0.32 397.695 69.945 ;
    RECT 396.495 0.32 397.125 69.945 ;
    RECT 394.945 0.32 396.145 69.945 ;
    RECT 394.365 0.32 394.595 69.945 ;
    RECT 393.395 0.32 394.015 69.945 ;
    RECT 392.415 0.32 393.045 69.945 ;
    RECT 391.845 0.32 392.065 69.945 ;
    RECT 391.275 0.32 391.495 69.945 ;
    RECT 390.295 0.32 390.925 69.945 ;
    RECT 388.745 0.32 389.945 69.945 ;
    RECT 388.165 0.32 388.395 69.945 ;
    RECT 387.195 0.32 387.815 69.945 ;
    RECT 386.215 0.32 386.845 69.945 ;
    RECT 385.645 0.32 385.865 69.945 ;
    RECT 385.075 0.32 385.295 69.945 ;
    RECT 384.095 0.32 384.725 69.945 ;
    RECT 382.545 0.32 383.745 69.945 ;
    RECT 381.965 0.32 382.195 69.945 ;
    RECT 380.995 0.32 381.615 69.945 ;
    RECT 380.015 0.32 380.645 69.945 ;
    RECT 379.445 0.32 379.665 69.945 ;
    RECT 378.875 0.32 379.095 69.945 ;
    RECT 377.895 0.32 378.525 69.945 ;
    RECT 376.345 0.32 377.545 69.945 ;
    RECT 375.765 0.32 375.995 69.945 ;
    RECT 374.795 0.32 375.415 69.945 ;
    RECT 373.815 0.32 374.445 69.945 ;
    RECT 373.245 0.32 373.465 69.945 ;
    RECT 372.675 0.32 372.895 69.945 ;
    RECT 371.695 0.32 372.325 69.945 ;
    RECT 370.145 0.32 371.345 69.945 ;
    RECT 369.565 0.32 369.795 69.945 ;
    RECT 368.595 0.32 369.215 69.945 ;
    RECT 367.615 0.32 368.245 69.945 ;
    RECT 367.045 0.32 367.265 69.945 ;
    RECT 366.475 0.32 366.695 69.945 ;
    RECT 365.495 0.32 366.125 69.945 ;
    RECT 363.945 0.32 365.145 69.945 ;
    RECT 363.365 0.32 363.595 69.945 ;
    RECT 362.395 0.32 363.015 69.945 ;
    RECT 361.415 0.32 362.045 69.945 ;
    RECT 360.845 0.32 361.065 69.945 ;
    RECT 360.275 0.32 360.495 69.945 ;
    RECT 359.295 0.32 359.925 69.945 ;
    RECT 357.745 0.32 358.945 69.945 ;
    RECT 357.165 0.32 357.395 69.945 ;
    RECT 356.195 0.32 356.815 69.945 ;
    RECT 355.215 0.32 355.845 69.945 ;
    RECT 354.645 0.32 354.865 69.945 ;
    RECT 354.075 0.32 354.295 69.945 ;
    RECT 353.095 0.32 353.725 69.945 ;
    RECT 351.545 0.32 352.745 69.945 ;
    RECT 350.965 0.32 351.195 69.945 ;
    RECT 349.995 0.32 350.615 69.945 ;
    RECT 349.015 0.32 349.645 69.945 ;
    RECT 348.445 0.32 348.665 69.945 ;
    RECT 347.875 0.32 348.095 69.945 ;
    RECT 346.895 0.32 347.525 69.945 ;
    RECT 345.345 0.32 346.545 69.945 ;
    RECT 344.765 0.32 344.995 69.945 ;
    RECT 343.795 0.32 344.415 69.945 ;
    RECT 342.815 0.32 343.445 69.945 ;
    RECT 342.245 0.32 342.465 69.945 ;
    RECT 341.675 0.32 341.895 69.945 ;
    RECT 340.695 0.32 341.325 69.945 ;
    RECT 339.145 0.32 340.345 69.945 ;
    RECT 338.565 0.32 338.795 69.945 ;
    RECT 337.595 0.32 338.215 69.945 ;
    RECT 336.615 0.32 337.245 69.945 ;
    RECT 336.045 0.32 336.265 69.945 ;
    RECT 335.475 0.32 335.695 69.945 ;
    RECT 334.495 0.32 335.125 69.945 ;
    RECT 332.945 0.32 334.145 69.945 ;
    RECT 332.365 0.32 332.595 69.945 ;
    RECT 331.395 0.32 332.015 69.945 ;
    RECT 330.415 0.32 331.045 69.945 ;
    RECT 329.845 0.32 330.065 69.945 ;
    RECT 329.275 0.32 329.495 69.945 ;
    RECT 328.295 0.32 328.925 69.945 ;
    RECT 326.745 0.32 327.945 69.945 ;
    RECT 326.165 0.32 326.395 69.945 ;
    RECT 325.195 0.32 325.815 69.945 ;
    RECT 324.215 0.32 324.845 69.945 ;
    RECT 323.645 0.32 323.865 69.945 ;
    RECT 323.075 0.32 323.295 69.945 ;
    RECT 322.095 0.32 322.725 69.945 ;
    RECT 320.545 0.32 321.745 69.945 ;
    RECT 319.965 0.32 320.195 69.945 ;
    RECT 318.995 0.32 319.615 69.945 ;
    RECT 318.015 0.32 318.645 69.945 ;
    RECT 317.445 0.32 317.665 69.945 ;
    RECT 316.875 0.32 317.095 69.945 ;
    RECT 315.895 0.32 316.525 69.945 ;
    RECT 314.345 0.32 315.545 69.945 ;
    RECT 313.765 0.32 313.995 69.945 ;
    RECT 312.795 0.32 313.415 69.945 ;
    RECT 311.815 0.32 312.445 69.945 ;
    RECT 311.245 0.32 311.465 69.945 ;
    RECT 310.675 0.32 310.895 69.945 ;
    RECT 309.695 0.32 310.325 69.945 ;
    RECT 308.145 0.32 309.345 69.945 ;
    RECT 307.565 0.32 307.795 69.945 ;
    RECT 306.595 0.32 307.215 69.945 ;
    RECT 305.615 0.32 306.245 69.945 ;
    RECT 305.045 0.32 305.265 69.945 ;
    RECT 304.475 0.32 304.695 69.945 ;
    RECT 303.495 0.32 304.125 69.945 ;
    RECT 301.945 0.32 303.145 69.945 ;
    RECT 301.365 0.32 301.595 69.945 ;
    RECT 300.395 0.32 301.015 69.945 ;
    RECT 299.415 0.32 300.045 69.945 ;
    RECT 298.845 0.32 299.065 69.945 ;
    RECT 298.275 0.32 298.495 69.945 ;
    RECT 297.295 0.32 297.925 69.945 ;
    RECT 295.745 0.32 296.945 69.945 ;
    RECT 295.165 0.32 295.395 69.945 ;
    RECT 294.195 0.32 294.815 69.945 ;
    RECT 293.215 0.32 293.845 69.945 ;
    RECT 292.645 0.32 292.865 69.945 ;
    RECT 292.075 0.32 292.295 69.945 ;
    RECT 291.095 0.32 291.725 69.945 ;
    RECT 289.545 0.32 290.745 69.945 ;
    RECT 288.965 0.32 289.195 69.945 ;
    RECT 287.995 0.32 288.615 69.945 ;
    RECT 287.015 0.32 287.645 69.945 ;
    RECT 286.445 0.32 286.665 69.945 ;
    RECT 285.875 0.32 286.095 69.945 ;
    RECT 284.895 0.32 285.525 69.945 ;
    RECT 283.345 0.32 284.545 69.945 ;
    RECT 282.765 0.32 282.995 69.945 ;
    RECT 281.795 0.32 282.415 69.945 ;
    RECT 280.815 0.32 281.445 69.945 ;
    RECT 280.245 0.32 280.465 69.945 ;
    RECT 279.675 0.32 279.895 69.945 ;
    RECT 278.695 0.32 279.325 69.945 ;
    RECT 277.145 0.32 278.345 69.945 ;
    RECT 276.565 0.32 276.795 69.945 ;
    RECT 275.595 0.32 276.215 69.945 ;
    RECT 274.615 0.32 275.245 69.945 ;
    RECT 274.045 0.32 274.265 69.945 ;
    RECT 273.475 0.32 273.695 69.945 ;
    RECT 272.495 0.32 273.125 69.945 ;
    RECT 270.945 0.32 272.145 69.945 ;
    RECT 270.365 0.32 270.595 69.945 ;
    RECT 269.395 0.32 270.015 69.945 ;
    RECT 268.415 0.32 269.045 69.945 ;
    RECT 267.845 0.32 268.065 69.945 ;
    RECT 267.275 0.32 267.495 69.945 ;
    RECT 266.295 0.32 266.925 69.945 ;
    RECT 264.745 0.32 265.945 69.945 ;
    RECT 264.165 0.32 264.395 69.945 ;
    RECT 263.195 0.32 263.815 69.945 ;
    RECT 262.215 0.32 262.845 69.945 ;
    RECT 261.645 0.32 261.865 69.945 ;
    RECT 261.075 0.32 261.295 69.945 ;
    RECT 260.095 0.32 260.725 69.945 ;
    RECT 258.545 0.32 259.745 69.945 ;
    RECT 257.965 0.32 258.195 69.945 ;
    RECT 256.995 0.32 257.615 69.945 ;
    RECT 256.015 0.32 256.645 69.945 ;
    RECT 255.445 0.32 255.665 69.945 ;
    RECT 254.875 0.32 255.095 69.945 ;
    RECT 253.895 0.32 254.525 69.945 ;
    RECT 252.345 0.32 253.545 69.945 ;
    RECT 251.765 0.32 251.995 69.945 ;
    RECT 250.795 0.32 251.415 69.945 ;
    RECT 249.815 0.32 250.445 69.945 ;
    RECT 249.245 0.32 249.465 69.945 ;
    RECT 248.675 0.32 248.895 69.945 ;
    RECT 247.695 0.32 248.325 69.945 ;
    RECT 246.145 0.32 247.345 69.945 ;
    RECT 245.565 0.32 245.795 69.945 ;
    RECT 244.595 0.32 245.215 69.945 ;
    RECT 243.615 0.32 244.245 69.945 ;
    RECT 243.045 0.32 243.265 69.945 ;
    RECT 241.305 0.32 242.695 69.945 ;
    RECT 240.515 0.32 240.955 69.945 ;
    RECT 239.515 0.32 240.165 69.945 ;
    RECT 235.96 0.32 236.82 69.945 ;
    RECT 235.4 0.32 235.48 69.945 ;
    RECT 233.84 0.32 234.27 69.945 ;
    RECT 232.705 0.32 233.49 69.945 ;
    RECT 231.44 0.32 232.225 69.945 ;
    RECT 230.675 0.32 230.98 69.945 ;
    RECT 229.505 0.32 229.935 69.945 ;
    RECT 227.565 0.32 227.995 69.945 ;
    RECT 226.915 0.32 227.215 69.945 ;
    RECT 225.32 0.32 225.79 69.945 ;
    RECT 224.52 0.32 224.97 69.945 ;
    RECT 223.95 0.32 224.17 69.945 ;
    RECT 222.29 0.32 223.49 69.945 ;
    RECT 221.78 0.32 221.94 69.945 ;
    RECT 221.0 0.32 221.43 69.945 ;
    RECT 220.49 0.32 220.65 69.945 ;
    RECT 218.94 0.32 220.14 69.945 ;
    RECT 218.26 0.32 218.48 69.945 ;
    RECT 217.46 0.32 217.91 69.945 ;
    RECT 216.64 0.32 217.11 69.945 ;
    RECT 215.215 0.32 215.515 69.945 ;
    RECT 214.435 0.32 214.865 69.945 ;
    RECT 212.495 0.32 212.925 69.945 ;
    RECT 211.45 0.32 211.755 69.945 ;
    RECT 210.205 0.32 210.99 69.945 ;
    RECT 208.94 0.32 209.725 69.945 ;
    RECT 208.16 0.32 208.59 69.945 ;
    RECT 206.95 0.32 207.03 69.945 ;
    RECT 205.61 0.32 206.47 69.945 ;
    RECT 202.265 0.32 202.915 69.945 ;
    RECT 201.475 0.32 201.915 69.945 ;
    RECT 199.735 0.32 201.125 69.945 ;
    RECT 199.165 0.32 199.385 69.945 ;
    RECT 198.185 0.32 198.815 69.945 ;
    RECT 197.215 0.32 197.835 69.945 ;
    RECT 196.635 0.32 196.865 69.945 ;
    RECT 195.085 0.32 196.285 69.945 ;
    RECT 194.105 0.32 194.735 69.945 ;
    RECT 193.535 0.32 193.755 69.945 ;
    RECT 192.965 0.32 193.185 69.945 ;
    RECT 191.985 0.32 192.615 69.945 ;
    RECT 191.015 0.32 191.635 69.945 ;
    RECT 190.435 0.32 190.665 69.945 ;
    RECT 188.885 0.32 190.085 69.945 ;
    RECT 187.905 0.32 188.535 69.945 ;
    RECT 187.335 0.32 187.555 69.945 ;
    RECT 186.765 0.32 186.985 69.945 ;
    RECT 185.785 0.32 186.415 69.945 ;
    RECT 184.815 0.32 185.435 69.945 ;
    RECT 184.235 0.32 184.465 69.945 ;
    RECT 182.685 0.32 183.885 69.945 ;
    RECT 181.705 0.32 182.335 69.945 ;
    RECT 181.135 0.32 181.355 69.945 ;
    RECT 180.565 0.32 180.785 69.945 ;
    RECT 179.585 0.32 180.215 69.945 ;
    RECT 178.615 0.32 179.235 69.945 ;
    RECT 178.035 0.32 178.265 69.945 ;
    RECT 176.485 0.32 177.685 69.945 ;
    RECT 175.505 0.32 176.135 69.945 ;
    RECT 174.935 0.32 175.155 69.945 ;
    RECT 174.365 0.32 174.585 69.945 ;
    RECT 173.385 0.32 174.015 69.945 ;
    RECT 172.415 0.32 173.035 69.945 ;
    RECT 171.835 0.32 172.065 69.945 ;
    RECT 170.285 0.32 171.485 69.945 ;
    RECT 169.305 0.32 169.935 69.945 ;
    RECT 168.735 0.32 168.955 69.945 ;
    RECT 168.165 0.32 168.385 69.945 ;
    RECT 167.185 0.32 167.815 69.945 ;
    RECT 166.215 0.32 166.835 69.945 ;
    RECT 165.635 0.32 165.865 69.945 ;
    RECT 164.085 0.32 165.285 69.945 ;
    RECT 163.105 0.32 163.735 69.945 ;
    RECT 162.535 0.32 162.755 69.945 ;
    RECT 161.965 0.32 162.185 69.945 ;
    RECT 160.985 0.32 161.615 69.945 ;
    RECT 160.015 0.32 160.635 69.945 ;
    RECT 159.435 0.32 159.665 69.945 ;
    RECT 157.885 0.32 159.085 69.945 ;
    RECT 156.905 0.32 157.535 69.945 ;
    RECT 156.335 0.32 156.555 69.945 ;
    RECT 155.765 0.32 155.985 69.945 ;
    RECT 154.785 0.32 155.415 69.945 ;
    RECT 153.815 0.32 154.435 69.945 ;
    RECT 153.235 0.32 153.465 69.945 ;
    RECT 151.685 0.32 152.885 69.945 ;
    RECT 150.705 0.32 151.335 69.945 ;
    RECT 150.135 0.32 150.355 69.945 ;
    RECT 149.565 0.32 149.785 69.945 ;
    RECT 148.585 0.32 149.215 69.945 ;
    RECT 147.615 0.32 148.235 69.945 ;
    RECT 147.035 0.32 147.265 69.945 ;
    RECT 145.485 0.32 146.685 69.945 ;
    RECT 144.505 0.32 145.135 69.945 ;
    RECT 143.935 0.32 144.155 69.945 ;
    RECT 143.365 0.32 143.585 69.945 ;
    RECT 142.385 0.32 143.015 69.945 ;
    RECT 141.415 0.32 142.035 69.945 ;
    RECT 140.835 0.32 141.065 69.945 ;
    RECT 139.285 0.32 140.485 69.945 ;
    RECT 138.305 0.32 138.935 69.945 ;
    RECT 137.735 0.32 137.955 69.945 ;
    RECT 137.165 0.32 137.385 69.945 ;
    RECT 136.185 0.32 136.815 69.945 ;
    RECT 135.215 0.32 135.835 69.945 ;
    RECT 134.635 0.32 134.865 69.945 ;
    RECT 133.085 0.32 134.285 69.945 ;
    RECT 132.105 0.32 132.735 69.945 ;
    RECT 131.535 0.32 131.755 69.945 ;
    RECT 130.965 0.32 131.185 69.945 ;
    RECT 129.985 0.32 130.615 69.945 ;
    RECT 129.015 0.32 129.635 69.945 ;
    RECT 128.435 0.32 128.665 69.945 ;
    RECT 126.885 0.32 128.085 69.945 ;
    RECT 125.905 0.32 126.535 69.945 ;
    RECT 125.335 0.32 125.555 69.945 ;
    RECT 124.765 0.32 124.985 69.945 ;
    RECT 123.785 0.32 124.415 69.945 ;
    RECT 122.815 0.32 123.435 69.945 ;
    RECT 122.235 0.32 122.465 69.945 ;
    RECT 120.685 0.32 121.885 69.945 ;
    RECT 119.705 0.32 120.335 69.945 ;
    RECT 119.135 0.32 119.355 69.945 ;
    RECT 118.565 0.32 118.785 69.945 ;
    RECT 117.585 0.32 118.215 69.945 ;
    RECT 116.615 0.32 117.235 69.945 ;
    RECT 116.035 0.32 116.265 69.945 ;
    RECT 114.485 0.32 115.685 69.945 ;
    RECT 113.505 0.32 114.135 69.945 ;
    RECT 112.935 0.32 113.155 69.945 ;
    RECT 112.365 0.32 112.585 69.945 ;
    RECT 111.385 0.32 112.015 69.945 ;
    RECT 110.415 0.32 111.035 69.945 ;
    RECT 109.835 0.32 110.065 69.945 ;
    RECT 108.285 0.32 109.485 69.945 ;
    RECT 107.305 0.32 107.935 69.945 ;
    RECT 106.735 0.32 106.955 69.945 ;
    RECT 106.165 0.32 106.385 69.945 ;
    RECT 105.185 0.32 105.815 69.945 ;
    RECT 104.215 0.32 104.835 69.945 ;
    RECT 103.635 0.32 103.865 69.945 ;
    RECT 102.085 0.32 103.285 69.945 ;
    RECT 101.105 0.32 101.735 69.945 ;
    RECT 100.535 0.32 100.755 69.945 ;
    RECT 99.965 0.32 100.185 69.945 ;
    RECT 98.985 0.32 99.615 69.945 ;
    RECT 98.015 0.32 98.635 69.945 ;
    RECT 97.435 0.32 97.665 69.945 ;
    RECT 95.885 0.32 97.085 69.945 ;
    RECT 94.905 0.32 95.535 69.945 ;
    RECT 94.335 0.32 94.555 69.945 ;
    RECT 93.765 0.32 93.985 69.945 ;
    RECT 92.785 0.32 93.415 69.945 ;
    RECT 91.815 0.32 92.435 69.945 ;
    RECT 91.235 0.32 91.465 69.945 ;
    RECT 89.685 0.32 90.885 69.945 ;
    RECT 88.705 0.32 89.335 69.945 ;
    RECT 88.135 0.32 88.355 69.945 ;
    RECT 87.565 0.32 87.785 69.945 ;
    RECT 86.585 0.32 87.215 69.945 ;
    RECT 85.615 0.32 86.235 69.945 ;
    RECT 85.035 0.32 85.265 69.945 ;
    RECT 83.485 0.32 84.685 69.945 ;
    RECT 82.505 0.32 83.135 69.945 ;
    RECT 81.935 0.32 82.155 69.945 ;
    RECT 81.365 0.32 81.585 69.945 ;
    RECT 80.385 0.32 81.015 69.945 ;
    RECT 79.415 0.32 80.035 69.945 ;
    RECT 78.835 0.32 79.065 69.945 ;
    RECT 77.285 0.32 78.485 69.945 ;
    RECT 76.305 0.32 76.935 69.945 ;
    RECT 75.735 0.32 75.955 69.945 ;
    RECT 75.165 0.32 75.385 69.945 ;
    RECT 74.185 0.32 74.815 69.945 ;
    RECT 73.215 0.32 73.835 69.945 ;
    RECT 72.635 0.32 72.865 69.945 ;
    RECT 71.085 0.32 72.285 69.945 ;
    RECT 70.105 0.32 70.735 69.945 ;
    RECT 69.535 0.32 69.755 69.945 ;
    RECT 68.965 0.32 69.185 69.945 ;
    RECT 67.985 0.32 68.615 69.945 ;
    RECT 67.015 0.32 67.635 69.945 ;
    RECT 66.435 0.32 66.665 69.945 ;
    RECT 64.885 0.32 66.085 69.945 ;
    RECT 63.905 0.32 64.535 69.945 ;
    RECT 63.335 0.32 63.555 69.945 ;
    RECT 62.765 0.32 62.985 69.945 ;
    RECT 61.785 0.32 62.415 69.945 ;
    RECT 60.815 0.32 61.435 69.945 ;
    RECT 60.235 0.32 60.465 69.945 ;
    RECT 58.685 0.32 59.885 69.945 ;
    RECT 57.705 0.32 58.335 69.945 ;
    RECT 57.135 0.32 57.355 69.945 ;
    RECT 56.565 0.32 56.785 69.945 ;
    RECT 55.585 0.32 56.215 69.945 ;
    RECT 54.615 0.32 55.235 69.945 ;
    RECT 54.035 0.32 54.265 69.945 ;
    RECT 52.485 0.32 53.685 69.945 ;
    RECT 51.505 0.32 52.135 69.945 ;
    RECT 50.935 0.32 51.155 69.945 ;
    RECT 50.365 0.32 50.585 69.945 ;
    RECT 49.385 0.32 50.015 69.945 ;
    RECT 48.415 0.32 49.035 69.945 ;
    RECT 47.835 0.32 48.065 69.945 ;
    RECT 46.285 0.32 47.485 69.945 ;
    RECT 45.305 0.32 45.935 69.945 ;
    RECT 44.735 0.32 44.955 69.945 ;
    RECT 44.165 0.32 44.385 69.945 ;
    RECT 43.185 0.32 43.815 69.945 ;
    RECT 42.215 0.32 42.835 69.945 ;
    RECT 41.635 0.32 41.865 69.945 ;
    RECT 40.085 0.32 41.285 69.945 ;
    RECT 39.105 0.32 39.735 69.945 ;
    RECT 38.535 0.32 38.755 69.945 ;
    RECT 37.965 0.32 38.185 69.945 ;
    RECT 36.985 0.32 37.615 69.945 ;
    RECT 36.015 0.32 36.635 69.945 ;
    RECT 35.435 0.32 35.665 69.945 ;
    RECT 33.885 0.32 35.085 69.945 ;
    RECT 32.905 0.32 33.535 69.945 ;
    RECT 32.335 0.32 32.555 69.945 ;
    RECT 31.765 0.32 31.985 69.945 ;
    RECT 30.785 0.32 31.415 69.945 ;
    RECT 29.815 0.32 30.435 69.945 ;
    RECT 29.235 0.32 29.465 69.945 ;
    RECT 27.685 0.32 28.885 69.945 ;
    RECT 26.705 0.32 27.335 69.945 ;
    RECT 26.135 0.32 26.355 69.945 ;
    RECT 25.565 0.32 25.785 69.945 ;
    RECT 24.585 0.32 25.215 69.945 ;
    RECT 23.615 0.32 24.235 69.945 ;
    RECT 23.035 0.32 23.265 69.945 ;
    RECT 21.485 0.32 22.685 69.945 ;
    RECT 20.505 0.32 21.135 69.945 ;
    RECT 19.935 0.32 20.155 69.945 ;
    RECT 19.365 0.32 19.585 69.945 ;
    RECT 18.385 0.32 19.015 69.945 ;
    RECT 17.415 0.32 18.035 69.945 ;
    RECT 16.835 0.32 17.065 69.945 ;
    RECT 15.285 0.32 16.485 69.945 ;
    RECT 14.305 0.32 14.935 69.945 ;
    RECT 13.735 0.32 13.955 69.945 ;
    RECT 13.165 0.32 13.385 69.945 ;
    RECT 12.185 0.32 12.815 69.945 ;
    RECT 11.215 0.32 11.835 69.945 ;
    RECT 10.635 0.32 10.865 69.945 ;
    RECT 9.085 0.32 10.285 69.945 ;
    RECT 8.105 0.32 8.735 69.945 ;
    RECT 7.535 0.32 7.755 69.945 ;
    RECT 6.965 0.32 7.185 69.945 ;
    RECT 5.985 0.32 6.615 69.945 ;
    RECT 5.015 0.32 5.635 69.945 ;
    RECT 4.435 0.32 4.665 69.945 ;
    RECT 2.885 0.32 4.085 69.945 ;
    RECT 1.905 0.32 2.535 69.945 ;
    RECT 1.335 0.32 1.555 69.945 ;
    RECT 0.0 0.32 0.985 69.945 ;
    END
  END SRAMdpw64d256

END LIBRARY

